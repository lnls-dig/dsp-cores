--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_1482f9e8df81448a.vhd when simulating
-- the core, addsb_11_0_1482f9e8df81448a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_1482f9e8df81448a IS
  PORT (
    a : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(26 DOWNTO 0)
  );
END addsb_11_0_1482f9e8df81448a;

ARCHITECTURE addsb_11_0_1482f9e8df81448a_a OF addsb_11_0_1482f9e8df81448a IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_1482f9e8df81448a
  PORT (
    a : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(26 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_1482f9e8df81448a USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 27,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000000000000",
      c_b_width => 27,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 27,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_1482f9e8df81448a
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_1482f9e8df81448a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_239e4f614ba09ab1.vhd when simulating
-- the core, addsb_11_0_239e4f614ba09ab1. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_239e4f614ba09ab1 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END addsb_11_0_239e4f614ba09ab1;

ARCHITECTURE addsb_11_0_239e4f614ba09ab1_a OF addsb_11_0_239e4f614ba09ab1 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_239e4f614ba09ab1
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_239e4f614ba09ab1 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 26,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000000000",
      c_b_width => 26,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 26,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_239e4f614ba09ab1
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_239e4f614ba09ab1_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_2f1626aeedb3c308.vhd when simulating
-- the core, addsb_11_0_2f1626aeedb3c308. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_2f1626aeedb3c308 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(26 DOWNTO 0)
  );
END addsb_11_0_2f1626aeedb3c308;

ARCHITECTURE addsb_11_0_2f1626aeedb3c308_a OF addsb_11_0_2f1626aeedb3c308 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_2f1626aeedb3c308
  PORT (
    a : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(26 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_2f1626aeedb3c308 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 27,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000000000000000000000",
      c_b_width => 27,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 27,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_2f1626aeedb3c308
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_2f1626aeedb3c308_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cc_cmplr_v3_0_2d327f6921329141.vhd when simulating
-- the core, cc_cmplr_v3_0_2d327f6921329141. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cc_cmplr_v3_0_2d327f6921329141 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC
  );
END cc_cmplr_v3_0_2d327f6921329141;

ARCHITECTURE cc_cmplr_v3_0_2d327f6921329141_a OF cc_cmplr_v3_0_2d327f6921329141 IS
-- synthesis translate_off
COMPONENT wrapped_cc_cmplr_v3_0_2d327f6921329141
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cc_cmplr_v3_0_2d327f6921329141 USE ENTITY XilinxCoreLib.cic_compiler_v3_0(behavioral)
    GENERIC MAP (
      c_c1 => 30,
      c_c2 => 29,
      c_c3 => 28,
      c_c4 => 27,
      c_c5 => 27,
      c_c6 => 0,
      c_clk_freq => 1,
      c_component_name => "cc_cmplr_v3_0_2d327f6921329141",
      c_diff_delay => 2,
      c_family => "virtex6",
      c_filter_type => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_dout_tready => 0,
      c_has_rounding => 0,
      c_i1 => 81,
      c_i2 => 69,
      c_i3 => 57,
      c_i4 => 46,
      c_i5 => 35,
      c_i6 => 0,
      c_input_width => 24,
      c_m_axis_data_tdata_width => 24,
      c_m_axis_data_tuser_width => 1,
      c_max_rate => 2500,
      c_min_rate => 2500,
      c_num_channels => 1,
      c_num_stages => 5,
      c_output_width => 24,
      c_rate => 2500,
      c_rate_type => 0,
      c_s_axis_config_tdata_width => 1,
      c_s_axis_data_tdata_width => 24,
      c_sample_freq => 1,
      c_use_dsp => 1,
      c_use_streaming_interface => 1,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cc_cmplr_v3_0_2d327f6921329141
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tdata => s_axis_data_tdata,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid
  );
-- synthesis translate_on

END cc_cmplr_v3_0_2d327f6921329141_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cc_cmplr_v3_0_75f3b28f5ac4aa5e.vhd when simulating
-- the core, cc_cmplr_v3_0_75f3b28f5ac4aa5e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cc_cmplr_v3_0_75f3b28f5ac4aa5e IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC
  );
END cc_cmplr_v3_0_75f3b28f5ac4aa5e;

ARCHITECTURE cc_cmplr_v3_0_75f3b28f5ac4aa5e_a OF cc_cmplr_v3_0_75f3b28f5ac4aa5e IS
-- synthesis translate_off
COMPONENT wrapped_cc_cmplr_v3_0_75f3b28f5ac4aa5e
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cc_cmplr_v3_0_75f3b28f5ac4aa5e USE ENTITY XilinxCoreLib.cic_compiler_v3_0(behavioral)
    GENERIC MAP (
      c_c1 => 31,
      c_c2 => 30,
      c_c3 => 29,
      c_c4 => 28,
      c_c5 => 28,
      c_c6 => 0,
      c_clk_freq => 1,
      c_component_name => "cc_cmplr_v3_0_75f3b28f5ac4aa5e",
      c_diff_delay => 2,
      c_family => "virtex6",
      c_filter_type => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_dout_tready => 0,
      c_has_rounding => 0,
      c_i1 => 77,
      c_i2 => 66,
      c_i3 => 55,
      c_i4 => 45,
      c_i5 => 36,
      c_i6 => 0,
      c_input_width => 24,
      c_m_axis_data_tdata_width => 32,
      c_m_axis_data_tuser_width => 1,
      c_max_rate => 1113,
      c_min_rate => 1113,
      c_num_channels => 1,
      c_num_stages => 5,
      c_output_width => 25,
      c_rate => 1113,
      c_rate_type => 0,
      c_s_axis_config_tdata_width => 1,
      c_s_axis_data_tdata_width => 24,
      c_sample_freq => 1,
      c_use_dsp => 1,
      c_use_streaming_interface => 1,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cc_cmplr_v3_0_75f3b28f5ac4aa5e
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tdata => s_axis_data_tdata,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid
  );
-- synthesis translate_on

END cc_cmplr_v3_0_75f3b28f5ac4aa5e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cmpy_v5_0_3b811ae68acefe54.vhd when simulating
-- the core, cmpy_v5_0_3b811ae68acefe54. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cmpy_v5_0_3b811ae68acefe54 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_a_tvalid : IN STD_LOGIC;
    s_axis_a_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    s_axis_b_tvalid : IN STD_LOGIC;
    s_axis_b_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END cmpy_v5_0_3b811ae68acefe54;

ARCHITECTURE cmpy_v5_0_3b811ae68acefe54_a OF cmpy_v5_0_3b811ae68acefe54 IS
-- synthesis translate_off
COMPONENT wrapped_cmpy_v5_0_3b811ae68acefe54
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_a_tvalid : IN STD_LOGIC;
    s_axis_a_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    s_axis_b_tvalid : IN STD_LOGIC;
    s_axis_b_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cmpy_v5_0_3b811ae68acefe54 USE ENTITY XilinxCoreLib.cmpy_v5_0(behavioral)
    GENERIC MAP (
      c_a_width => 24,
      c_b_width => 24,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_s_axis_a_tlast => 0,
      c_has_s_axis_a_tuser => 0,
      c_has_s_axis_b_tlast => 0,
      c_has_s_axis_b_tuser => 0,
      c_has_s_axis_ctrl_tlast => 0,
      c_has_s_axis_ctrl_tuser => 0,
      c_latency => 6,
      c_m_axis_dout_tdata_width => 48,
      c_m_axis_dout_tuser_width => 1,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_width => 24,
      c_s_axis_a_tdata_width => 48,
      c_s_axis_a_tuser_width => 1,
      c_s_axis_b_tdata_width => 48,
      c_s_axis_b_tuser_width => 1,
      c_s_axis_ctrl_tdata_width => 8,
      c_s_axis_ctrl_tuser_width => 1,
      c_throttle_scheme => 3,
      c_tlast_resolution => 0,
      c_verbosity => 0,
      c_xdevice => "xc6vlx240t",
      c_xdevicefamily => "virtex6",
      has_negate => 0,
      round => 0,
      single_output => 0,
      use_dsp_cascades => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cmpy_v5_0_3b811ae68acefe54
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_a_tvalid => s_axis_a_tvalid,
    s_axis_a_tdata => s_axis_a_tdata,
    s_axis_b_tvalid => s_axis_b_tvalid,
    s_axis_b_tdata => s_axis_b_tdata,
    m_axis_dout_tvalid => m_axis_dout_tvalid,
    m_axis_dout_tdata => m_axis_dout_tdata
  );
-- synthesis translate_on

END cmpy_v5_0_3b811ae68acefe54_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file crdc_v5_0_ac582be577bf89c0.vhd when simulating
-- the core, crdc_v5_0_ac582be577bf89c0. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY crdc_v5_0_ac582be577bf89c0 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_cartesian_tvalid : IN STD_LOGIC;
    s_axis_cartesian_tdata : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
  );
END crdc_v5_0_ac582be577bf89c0;

ARCHITECTURE crdc_v5_0_ac582be577bf89c0_a OF crdc_v5_0_ac582be577bf89c0 IS
-- synthesis translate_off
COMPONENT wrapped_crdc_v5_0_ac582be577bf89c0
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_cartesian_tvalid : IN STD_LOGIC;
    s_axis_cartesian_tdata : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_crdc_v5_0_ac582be577bf89c0 USE ENTITY XilinxCoreLib.cordic_v5_0(behavioral)
    GENERIC MAP (
      c_architecture => 2,
      c_coarse_rotate => 1,
      c_cordic_function => 1,
      c_data_format => 0,
      c_has_aclk => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_s_axis_cartesian => 1,
      c_has_s_axis_cartesian_tlast => 0,
      c_has_s_axis_cartesian_tuser => 0,
      c_has_s_axis_phase => 0,
      c_has_s_axis_phase_tlast => 0,
      c_has_s_axis_phase_tuser => 0,
      c_input_width => 25,
      c_iterations => 0,
      c_m_axis_dout_tdata_width => 64,
      c_m_axis_dout_tuser_width => 1,
      c_output_width => 25,
      c_phase_format => 0,
      c_pipeline_mode => -2,
      c_precision => 0,
      c_round_mode => 3,
      c_s_axis_cartesian_tdata_width => 64,
      c_s_axis_cartesian_tuser_width => 1,
      c_s_axis_phase_tdata_width => 32,
      c_s_axis_phase_tuser_width => 1,
      c_scale_comp => 2,
      c_throttle_scheme => 3,
      c_tlast_resolution => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_crdc_v5_0_ac582be577bf89c0
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_cartesian_tvalid => s_axis_cartesian_tvalid,
    s_axis_cartesian_tdata => s_axis_cartesian_tdata,
    m_axis_dout_tvalid => m_axis_dout_tvalid,
    m_axis_dout_tdata => m_axis_dout_tdata
  );
-- synthesis translate_on

END crdc_v5_0_ac582be577bf89c0_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dds_cmplr_v5_0_61b575ede3cdcc97.vhd when simulating
-- the core, dds_cmplr_v5_0_61b575ede3cdcc97. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dds_cmplr_v5_0_61b575ede3cdcc97 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tready : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END dds_cmplr_v5_0_61b575ede3cdcc97;

ARCHITECTURE dds_cmplr_v5_0_61b575ede3cdcc97_a OF dds_cmplr_v5_0_61b575ede3cdcc97 IS
-- synthesis translate_off
COMPONENT wrapped_dds_cmplr_v5_0_61b575ede3cdcc97
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tready : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dds_cmplr_v5_0_61b575ede3cdcc97 USE ENTITY XilinxCoreLib.dds_compiler_v5_0(behavioral)
    GENERIC MAP (
      c_accumulator_width => 30,
      c_amplitude => 1,
      c_chan_width => 1,
      c_channels => 1,
      c_debug_interface => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_channel_index => 0,
      c_has_m_data => 1,
      c_has_m_phase => 0,
      c_has_phase_out => 0,
      c_has_phasegen => 1,
      c_has_s_config => 0,
      c_has_s_phase => 0,
      c_has_sincos => 1,
      c_has_tlast => 0,
      c_has_tready => 1,
      c_latency => 12,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 48,
      c_m_data_tuser_width => 1,
      c_m_phase_has_tuser => 0,
      c_m_phase_tdata_width => 1,
      c_m_phase_tuser_width => 1,
      c_mem_type => 1,
      c_negative_cosine => 0,
      c_negative_sine => 1,
      c_noise_shaping => 2,
      c_optimise_goal => 0,
      c_output_width => 24,
      c_outputs_required => 2,
      c_phase_angle_width => 11,
      c_phase_increment => 2,
      c_phase_increment_value => "1110101000001110101000001110,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0",
      c_phase_offset => 2,
      c_phase_offset_value => "0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0",
      c_por_mode => 0,
      c_s_config_sync_mode => 0,
      c_s_config_tdata_width => 1,
      c_s_phase_has_tuser => 0,
      c_s_phase_tdata_width => 1,
      c_s_phase_tuser_width => 1,
      c_use_dsp48 => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dds_cmplr_v5_0_61b575ede3cdcc97
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tready => m_axis_data_tready,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END dds_cmplr_v5_0_61b575ede3cdcc97_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.87xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v4_0_5ce7b020ea0b7ee9.vhd
-- /___/   /\     Timestamp: Tue Mar 26 15:36:14 2013
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -w -sim -ofmt vhdl C:/TEMP/sysgentmp-lucas.russo/cg_wk/c7a65db6ef26e2610/tmp/_cg/dv_gn_v4_0_5ce7b020ea0b7ee9.ngc C:/TEMP/sysgentmp-lucas.russo/cg_wk/c7a65db6ef26e2610/tmp/_cg/dv_gn_v4_0_5ce7b020ea0b7ee9.vhd 
-- Device	: 6vlx240tff1156-1
-- Input file	: C:/TEMP/sysgentmp-lucas.russo/cg_wk/c7a65db6ef26e2610/tmp/_cg/dv_gn_v4_0_5ce7b020ea0b7ee9.ngc
-- Output file	: C:/TEMP/sysgentmp-lucas.russo/cg_wk/c7a65db6ef26e2610/tmp/_cg/dv_gn_v4_0_5ce7b020ea0b7ee9.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v4_0_5ce7b020ea0b7ee9
-- Xilinx	: c:\xilinx\13.4\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v4_0_5ce7b020ea0b7ee9 is
  port (
    aclk : in STD_LOGIC := 'X'; 
    aclken : in STD_LOGIC := 'X'; 
    s_axis_divisor_tvalid : in STD_LOGIC := 'X'; 
    s_axis_dividend_tvalid : in STD_LOGIC := 'X'; 
    s_axis_divisor_tready : out STD_LOGIC; 
    s_axis_dividend_tready : out STD_LOGIC; 
    m_axis_dout_tvalid : out STD_LOGIC; 
    s_axis_divisor_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    s_axis_dividend_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    m_axis_dout_tdata : out STD_LOGIC_VECTOR ( 79 downto 0 ) 
  );
end dv_gn_v4_0_5ce7b020ea0b7ee9;

architecture STRUCTURE of dv_gn_v4_0_5ce7b020ea0b7ee9 is
  signal NlwRenamedSig_OI_s_axis_dividend_tready : STD_LOGIC; 
  signal N0 : STD_LOGIC; 
  signal U0_i_synth_valid_access_in : STD_LOGIC; 
  signal U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_39_135 : STD_LOGIC; 
  signal U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_first_q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_BYPASS_INV_403_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_BYPASS_INV_400_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_carrycascout : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_negate_balance_opt_has_pipe_first_q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_bypass_balance_opt_has_pipe_first_q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_pipe_4_418 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_last_digit_518 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_28_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_29_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_30_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_31_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_32_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_33_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_34_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_35_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_36_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_37_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_38_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_39_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_40_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_41_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_42_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_43_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_44_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_45_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_46_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_47_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_48_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_49_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_50_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_51_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_pipe_10_688 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_bdd0 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_A_Z_DET_RTL_delay_0_0_893 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_a : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_b : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_int : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_op_a : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_int_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_all_bits_zero_del : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_OP_DEL_RTL_delay_0_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_carry_rnd2 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_round_rnd1 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_0_GND_233_o_MUX_252_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_1_GND_233_o_MUX_251_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_2_GND_233_o_MUX_250_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_3_GND_233_o_MUX_249_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_4_GND_233_o_MUX_248_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_5_GND_233_o_MUX_247_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_6_GND_233_o_MUX_246_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_7_GND_233_o_MUX_245_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_8_GND_233_o_MUX_244_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_9_GND_233_o_MUX_243_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_10_GND_233_o_MUX_242_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_11_GND_233_o_MUX_241_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_12_GND_233_o_MUX_240_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_13_GND_233_o_MUX_239_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_14_GND_233_o_MUX_238_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_15_GND_233_o_MUX_237_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_16_GND_233_o_MUX_236_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_17_GND_233_o_MUX_235_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_18_GND_233_o_MUX_234_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_19_GND_233_o_MUX_233_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_20_GND_233_o_MUX_232_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_21_GND_233_o_MUX_231_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_22_GND_233_o_MUX_230_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_23_GND_233_o_MUX_229_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_24_GND_233_o_MUX_228_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_25_GND_233_o_MUX_177_o : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_first_q_1227 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_div_by_zero_del_opt_has_pipe_first_q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_33_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_34_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_35_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_36_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_37_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_38_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_39_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_40_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_41_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_42_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_43_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_44_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_45_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_46_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_47_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_48_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_49_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_50_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_51_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_52_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_53_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_54_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_55_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_56_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_57_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_58_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_59_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_60_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_61_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_62_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_63_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_64_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_65_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_66_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_67_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_68_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_69_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_70_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_71_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_72_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_73_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_74_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_75_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_76_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_77_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_78_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_79_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_80_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_81_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_82_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_83_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_84_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_85_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_86_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_87_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_88_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_33_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_34_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_35_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_36_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_37_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_38_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_39_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_40_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_53_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_54_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_55_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_56_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_57_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_58_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_59_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_60_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_61_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_62_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_63_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_64_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_65_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_66_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_67_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_68_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_69_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_70_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_71_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_72_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_73_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_74_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_75_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_76_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_77_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_78_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_79_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_80_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_81_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_82_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_83_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_84_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_85_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_86_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_87_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_88_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_89_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_first_q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_subtract_reg_opt_has_pipe_first_q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_33_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_34_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_35_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_36_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_37_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_38_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_39_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_40_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_41_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_42_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_43_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_44_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_45_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_46_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_47_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_33_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_47_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_19_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_20_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_21_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_22_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_23_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_24_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_25_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_26_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_27_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_28_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_29_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_30_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_31_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_32_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_17_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_18_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_0_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_1_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_2_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_3_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_4_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_5_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_14_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_15_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_1_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_2_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_3_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_4_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_5_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_6_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_7_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_8_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_9_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_10_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_11_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_12_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_13_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_14_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_15_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_16_Q : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_7_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_8_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_9_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_10_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_11_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_12_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_13_Q : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX_rt_2543 : STD_LOGIC;
 
  signal U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0_2544 : STD_LOGIC; 
  signal U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1_2545 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4_2546 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26_2547 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25_2548 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22_2549 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24_2550 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23_2551 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19_2552 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21_2553 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20_2554 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16_2555 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18_2556 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17_2557 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15_2558 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14_2559 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13_2560 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12_2561 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9_2562 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11_2563 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10_2564 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6_2565 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8_2566 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7_2567 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3_2568 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5_2569 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4_2570 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2_2571 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1_2572 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0_2573 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1_2574 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20_2575 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0_2576 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1_2577 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q_2578 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15_2579 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14_2580 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16_2581 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15_2582 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13_2583 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12_2584 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11_2585 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10_2586 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7_2587 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9_2588 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8_2589 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4_2590 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6_2591 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5_2592 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1_2593 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3_2594 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2_2595 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0_2596 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26_2597 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25_2598 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24_2599 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21_2600 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23_2601 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22_2602 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18_2603 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20_2604 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19_2605 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17_2606 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16_2607 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5_2608 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4_2609 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1_2610 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3_2611 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2_2612 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1_2613 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0_2614 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3_2615 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12_2616 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13_2617 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9_2618 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11_2619 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10_2620 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6_2621 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8_2622 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7_2623 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16_2624 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18_2625 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17_2626 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15_2627 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14_2628 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13_2629 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12_2630 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9_2631 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11_2632 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10_2633 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6_2634 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8_2635 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7_2636 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3_2637 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5_2638 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4_2639 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2_2640 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1_2641 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0_2642 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2643 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2644 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2645 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2646 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2647 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2648 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2649 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2650 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2651 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2652 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2653 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2654 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2655 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2656 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2657 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2658 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2659 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2660 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2661 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2662 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2663 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2664 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2665 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2666 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2667 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2668 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2669 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2670 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2671 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2672 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2673 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2674 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2675 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2676 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2677 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2678 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2679 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2680 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2681 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2682 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2683 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2684 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2685 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2686 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2687 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2688 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2689 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2690 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37_2691 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36_2692 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35_2693 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34_2694 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31_2695 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33_2696 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32_2697 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28_2698 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30_2699 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29_2700 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25_2701 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27_2702 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26_2703 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24_2704 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23_2705 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22_2706 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21_2707 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18_2708 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20_2709 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19_2710 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15_2711 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17_2712 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16_2713 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12_2714 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14_2715 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13_2716 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9_2717 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11_2718 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10_2719 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6_2720 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8_2721 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7_2722 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3_2723 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5_2724 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4_2725 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0_2726 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2_2727 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1_2728 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10_2729 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15_2730 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14_2731 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13_2732 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12_2733 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11_2734 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8_2735 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10_2736 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9_2737 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5_2738 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7_2739 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6_2740 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2_2741 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4_2742 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3_2743 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1_2744 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0_2745 : STD_LOGIC; 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2_2746 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3_2747 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4_2748 : STD_LOGIC;
 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit_2749 : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_27_NO_RLOCS_Q_XOR_SUM_XOR_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_1_MUX_OP_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_2_MUX_OP_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP_O_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_CASCADEOUTA_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_CASCADEOUTB_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPA_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPA_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPB_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPB_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4_Q15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED : STD_LOGIC;
 
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED : STD_LOGIC;
 
  signal NlwRenamedSignal_m_axis_dout_tdata : STD_LOGIC_VECTOR ( 72 downto 72 ); 
  signal NlwRenamedSig_OI_m_axis_dout_tdata : STD_LOGIC_VECTOR ( 59 downto 36 ); 
  signal NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 47 downto 12 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout : STD_LOGIC_VECTOR3 ( 0 downto 0 , 0 downto 0 , 29 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi : STD_LOGIC_VECTOR3 ( 0 downto 0 , 0 downto 0 , 16 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout : STD_LOGIC_VECTOR3 ( 0 downto 0 , 0 downto 0 , 47 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1 : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2 : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d : STD_LOGIC_VECTOR ( 37 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 11 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb : STD_LOGIC_VECTOR ( 33 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2 : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout1 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout2 : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset : STD_LOGIC_VECTOR ( 16 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d : STD_LOGIC_VECTOR ( 21 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_pre_del_offset : STD_LOGIC_VECTOR ( 16 downto 16 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line : STD_LOGIC_VECTOR ( 12 downto 2 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 4 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit : STD_LOGIC_VECTOR ( 15 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom : STD_LOGIC_VECTOR ( 27 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d : STD_LOGIC_VECTOR ( 18 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d : STD_LOGIC_VECTOR ( 26 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate : STD_LOGIC_VECTOR ( 18 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op : STD_LOGIC_VECTOR ( 25 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9 : STD_LOGIC_VECTOR ( 26 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Madd_EXP_OUT_lut : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0 : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0 : STD_LOGIC_VECTOR ( 12 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0 : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0 : STD_LOGIC_VECTOR ( 26 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0 : STD_LOGIC_VECTOR ( 26 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a : STD_LOGIC_VECTOR ( 25 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp : STD_LOGIC_VECTOR ( 5 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int : STD_LOGIC_VECTOR ( 26 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry : STD_LOGIC_VECTOR ( 27 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry : STD_LOGIC_VECTOR ( 8 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry : STD_LOGIC_VECTOR ( 6 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_a_ip : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_carry : STD_LOGIC_VECTOR ( 2 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2 : STD_LOGIC_VECTOR ( 12 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1 : STD_LOGIC_VECTOR ( 12 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int : STD_LOGIC_VECTOR ( 12 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry : STD_LOGIC_VECTOR ( 12 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry : STD_LOGIC_VECTOR ( 13 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel : STD_LOGIC_VECTOR2 ( 0 downto 0 , 6 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux : STD_LOGIC_VECTOR ( 14 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave : STD_LOGIC_VECTOR2 ( 2 downto 0 , 18 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom : STD_LOGIC_VECTOR2 ( 2 downto 0 , 16 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom : STD_LOGIC_VECTOR2 ( 2 downto 0 , 15 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate : STD_LOGIC_VECTOR ( 17 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux : STD_LOGIC_VECTOR ( 17 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc : STD_LOGIC_VECTOR2 ( 2 downto 0 , 47 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave : STD_LOGIC_VECTOR2 ( 2 downto 0 , 18 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d : STD_LOGIC_VECTOR ( 29 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed : STD_LOGIC_VECTOR ( 33 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc : STD_LOGIC_VECTOR ( 47 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d : STD_LOGIC_VECTOR ( 17 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3 : STD_LOGIC_VECTOR ( 18 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d : STD_LOGIC_VECTOR ( 18 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op : STD_LOGIC_VECTOR2 ( 2 downto 2 , 15 downto 2 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op : STD_LOGIC_VECTOR ( 14 downto 1 ); 
  signal U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux : STD_LOGIC_VECTOR ( 18 downto 0 ); 
begin
  m_axis_dout_tdata(79) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(78) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(77) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(76) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(75) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(74) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(73) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(72) <= NlwRenamedSignal_m_axis_dout_tdata(72);
  m_axis_dout_tdata(59) <= NlwRenamedSig_OI_m_axis_dout_tdata(59);
  m_axis_dout_tdata(58) <= NlwRenamedSig_OI_m_axis_dout_tdata(58);
  m_axis_dout_tdata(57) <= NlwRenamedSig_OI_m_axis_dout_tdata(57);
  m_axis_dout_tdata(56) <= NlwRenamedSig_OI_m_axis_dout_tdata(56);
  m_axis_dout_tdata(55) <= NlwRenamedSig_OI_m_axis_dout_tdata(55);
  m_axis_dout_tdata(54) <= NlwRenamedSig_OI_m_axis_dout_tdata(54);
  m_axis_dout_tdata(53) <= NlwRenamedSig_OI_m_axis_dout_tdata(53);
  m_axis_dout_tdata(52) <= NlwRenamedSig_OI_m_axis_dout_tdata(52);
  m_axis_dout_tdata(51) <= NlwRenamedSig_OI_m_axis_dout_tdata(51);
  m_axis_dout_tdata(50) <= NlwRenamedSig_OI_m_axis_dout_tdata(50);
  m_axis_dout_tdata(49) <= NlwRenamedSig_OI_m_axis_dout_tdata(49);
  m_axis_dout_tdata(48) <= NlwRenamedSig_OI_m_axis_dout_tdata(48);
  m_axis_dout_tdata(47) <= NlwRenamedSig_OI_m_axis_dout_tdata(47);
  m_axis_dout_tdata(46) <= NlwRenamedSig_OI_m_axis_dout_tdata(46);
  m_axis_dout_tdata(45) <= NlwRenamedSig_OI_m_axis_dout_tdata(45);
  m_axis_dout_tdata(44) <= NlwRenamedSig_OI_m_axis_dout_tdata(44);
  m_axis_dout_tdata(43) <= NlwRenamedSig_OI_m_axis_dout_tdata(43);
  m_axis_dout_tdata(42) <= NlwRenamedSig_OI_m_axis_dout_tdata(42);
  m_axis_dout_tdata(41) <= NlwRenamedSig_OI_m_axis_dout_tdata(41);
  m_axis_dout_tdata(40) <= NlwRenamedSig_OI_m_axis_dout_tdata(40);
  m_axis_dout_tdata(39) <= NlwRenamedSig_OI_m_axis_dout_tdata(39);
  m_axis_dout_tdata(38) <= NlwRenamedSig_OI_m_axis_dout_tdata(38);
  m_axis_dout_tdata(37) <= NlwRenamedSig_OI_m_axis_dout_tdata(37);
  m_axis_dout_tdata(36) <= NlwRenamedSig_OI_m_axis_dout_tdata(36);
  m_axis_dout_tdata(35) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(47);
  m_axis_dout_tdata(34) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(46);
  m_axis_dout_tdata(33) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(45);
  m_axis_dout_tdata(32) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(44);
  m_axis_dout_tdata(31) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(43);
  m_axis_dout_tdata(30) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(42);
  m_axis_dout_tdata(29) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(41);
  m_axis_dout_tdata(28) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(40);
  m_axis_dout_tdata(27) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(39);
  m_axis_dout_tdata(26) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(38);
  m_axis_dout_tdata(25) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(37);
  m_axis_dout_tdata(24) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(36);
  m_axis_dout_tdata(23) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(35);
  m_axis_dout_tdata(22) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(34);
  m_axis_dout_tdata(21) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(33);
  m_axis_dout_tdata(20) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(32);
  m_axis_dout_tdata(19) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(31);
  m_axis_dout_tdata(18) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(30);
  m_axis_dout_tdata(17) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(29);
  m_axis_dout_tdata(16) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(28);
  m_axis_dout_tdata(15) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(27);
  m_axis_dout_tdata(14) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(26);
  m_axis_dout_tdata(13) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(25);
  m_axis_dout_tdata(12) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(24);
  m_axis_dout_tdata(11) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(23);
  m_axis_dout_tdata(10) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(22);
  m_axis_dout_tdata(9) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(21);
  m_axis_dout_tdata(8) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(20);
  m_axis_dout_tdata(7) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(19);
  m_axis_dout_tdata(6) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(18);
  m_axis_dout_tdata(5) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(17);
  m_axis_dout_tdata(4) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(16);
  m_axis_dout_tdata(3) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(15);
  m_axis_dout_tdata(2) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(14);
  m_axis_dout_tdata(1) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(13);
  m_axis_dout_tdata(0) <= 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(12);
  s_axis_divisor_tready <= NlwRenamedSig_OI_s_axis_dividend_tready;
  s_axis_dividend_tready <= NlwRenamedSig_OI_s_axis_dividend_tready;
  XST_VCC : VCC
    port map (
      P => N0
    );
  XST_GND : GND
    port map (
      G => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_valid_access_in,
      Q => U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1 : 
DSP48E1
    generic map(
      ACASCREG => 1,
      ADREG => 0,
      ALUMODEREG => 0,
      AREG => 1,
      AUTORESET_PATDET => "NO_RESET",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      DREG => 0,
      INMODEREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      USE_DPORT => FALSE,
      USE_MULT => "MULTIPLY",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEAD => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_MULTSIGNOUT_UNCONNECTED
,
      CEC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CED => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTD => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEA2 => aclken,
      CLK => aclk,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEM => aclken,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTINMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEINMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACOUT(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 29),
      ACOUT(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 28),
      ACOUT(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 27),
      ACOUT(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 26),
      ACOUT(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 25),
      ACOUT(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 24),
      ACOUT(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 23),
      ACOUT(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 22),
      ACOUT(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 21),
      ACOUT(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 20),
      ACOUT(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 19),
      ACOUT(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 18),
      ACOUT(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 17),
      ACOUT(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 16),
      ACOUT(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 15),
      ACOUT(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 14),
      ACOUT(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 13),
      ACOUT(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 12),
      ACOUT(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 11),
      ACOUT(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 10),
      ACOUT(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 9),
      ACOUT(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 8),
      ACOUT(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 7),
      ACOUT(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 6),
      ACOUT(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 5),
      ACOUT(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 4),
      ACOUT(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 3),
      ACOUT(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 2),
      ACOUT(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 1),
      ACOUT(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 0),
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_CARRYOUT_0_UNCONNECTED
,
      INMODE(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(16),
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(15),
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(14),
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(13),
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(12),
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(11),
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(10),
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(9),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(8),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(7),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(6),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(5),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(4),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(3),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(2),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(1),
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(0),
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_BCOUT_0_UNCONNECTED
,
      D(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_use_dsp48e1_iDSP48E1_P_17_UNCONNECTED
,
      P(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 16),
      P(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 15),
      P(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 14),
      P(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 13),
      P(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 12),
      P(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 11),
      P(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 10),
      P(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 9),
      P(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 8),
      P(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 7),
      P(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 6),
      P(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 5),
      P(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 4),
      P(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 3),
      P(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 2),
      P(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 1),
      P(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 0),
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(17),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(16),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(15),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(14),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(13),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(12),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(11),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(10),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(9),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(8),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(7),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(6),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(5),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(4),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(3),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(2),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(1),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(0),
      PCOUT(47) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 47),
      PCOUT(46) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 46),
      PCOUT(45) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 45),
      PCOUT(44) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 44),
      PCOUT(43) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 43),
      PCOUT(42) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 42),
      PCOUT(41) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 41),
      PCOUT(40) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 40),
      PCOUT(39) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 39),
      PCOUT(38) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 38),
      PCOUT(37) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 37),
      PCOUT(36) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 36),
      PCOUT(35) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 35),
      PCOUT(34) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 34),
      PCOUT(33) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 33),
      PCOUT(32) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 32),
      PCOUT(31) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 31),
      PCOUT(30) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 30),
      PCOUT(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 29),
      PCOUT(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 28),
      PCOUT(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 27),
      PCOUT(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 26),
      PCOUT(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 25),
      PCOUT(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 24),
      PCOUT(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 23),
      PCOUT(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 22),
      PCOUT(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 21),
      PCOUT(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 20),
      PCOUT(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 19),
      PCOUT(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 18),
      PCOUT(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 17),
      PCOUT(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 16),
      PCOUT(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 15),
      PCOUT(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 14),
      PCOUT(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 13),
      PCOUT(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 12),
      PCOUT(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 11),
      PCOUT(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 10),
      PCOUT(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 9),
      PCOUT(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 8),
      PCOUT(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 7),
      PCOUT(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 6),
      PCOUT(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 5),
      PCOUT(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 4),
      PCOUT(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 3),
      PCOUT(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 2),
      PCOUT(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 1),
      PCOUT(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 0),
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1 : 
DSP48E1
    generic map(
      ACASCREG => 1,
      ADREG => 0,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATDET => "NO_RESET",
      A_INPUT => "CASCADE",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      DREG => 0,
      INMODEREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      USE_DPORT => FALSE,
      USE_MULT => "MULTIPLY",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => aclken,
      CEAD => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_MULTSIGNOUT_UNCONNECTED
,
      CEC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CED => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTD => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CLK => aclk,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEM => aclken,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTINMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEINMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_ACOUT_0_UNCONNECTED
,
      OPMODE(6) => N0,
      OPMODE(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 47),
      PCIN(46) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 46),
      PCIN(45) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 45),
      PCIN(44) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 44),
      PCIN(43) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 43),
      PCIN(42) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 42),
      PCIN(41) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 41),
      PCIN(40) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 40),
      PCIN(39) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 39),
      PCIN(38) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 38),
      PCIN(37) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 37),
      PCIN(36) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 36),
      PCIN(35) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 35),
      PCIN(34) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 34),
      PCIN(33) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 33),
      PCIN(32) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 32),
      PCIN(31) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 31),
      PCIN(30) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 30),
      PCIN(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 29),
      PCIN(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 28),
      PCIN(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 27),
      PCIN(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 26),
      PCIN(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 25),
      PCIN(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 24),
      PCIN(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 23),
      PCIN(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 22),
      PCIN(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 21),
      PCIN(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 20),
      PCIN(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 19),
      PCIN(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 18),
      PCIN(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 17),
      PCIN(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 16),
      PCIN(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 15),
      PCIN(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 14),
      PCIN(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 13),
      PCIN(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 12),
      PCIN(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 11),
      PCIN(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 10),
      PCIN(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 9),
      PCIN(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 8),
      PCIN(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 7),
      PCIN(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 6),
      PCIN(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 5),
      PCIN(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 4),
      PCIN(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 3),
      PCIN(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 2),
      PCIN(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 1),
      PCIN(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pcout(0, 0, 0),
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_CARRYOUT_0_UNCONNECTED
,
      INMODE(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      INMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(26),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(25),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(24),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(23),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(22),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(21),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(20),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(19),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(18),
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(17),
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_BCOUT_0_UNCONNECTED
,
      D(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      D(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_P_11_UNCONNECTED
,
      P(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(27),
      P(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(26),
      P(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(25),
      P(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(24),
      P(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(23),
      P(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(22),
      P(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(21),
      P(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(20),
      P(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(19),
      P(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(18),
      P(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(17),
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_1_use_dsp48e1_iDSP48E1_PCOUT_0_UNCONNECTED
,
      ACIN(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 29),
      ACIN(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 28),
      ACIN(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 27),
      ACIN(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 26),
      ACIN(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 25),
      ACIN(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 24),
      ACIN(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 23),
      ACIN(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 22),
      ACIN(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 21),
      ACIN(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 20),
      ACIN(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 19),
      ACIN(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 18),
      ACIN(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 17),
      ACIN(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 16),
      ACIN(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 15),
      ACIN(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 14),
      ACIN(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 13),
      ACIN(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 12),
      ACIN(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 11),
      ACIN(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 10),
      ACIN(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 9),
      ACIN(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 8),
      ACIN(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 7),
      ACIN(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 6),
      ACIN(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 5),
      ACIN(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 4),
      ACIN(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 3),
      ACIN(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 2),
      ACIN(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 1),
      ACIN(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_acout(0, 0, 0),
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_bypass_balance_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_bypass_balance_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_negate_balance_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_negate_balance_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_10_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_9_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_8_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_7_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_6_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_5_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_4_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_3_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_10 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_2_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_11 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_1_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_12 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_0_Q
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_27_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(27)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_27_NO_RLOCS_Q_XOR_SUM_XOR_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_26_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(26)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_26_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(26)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(27)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_25_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(25)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(25),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_25_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(25)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(25),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_24_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(24)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(24),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_24_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(24)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(24),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_23_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(23)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(23),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_23_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(23)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(23),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_22_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(22)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(22),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_22_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(22)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(22),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_21_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(21)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(21),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_21_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(21)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(21),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_20_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(20)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(20),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_20_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(20)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(20),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_19_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(19)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(19),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_19_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(19)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(19),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_18_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(18)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(18),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_18_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(18)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(18),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_17_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(17)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(17),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_17_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(17)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(17),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_16_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(16)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(16),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_16_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(16)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(16),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_15_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(15)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(15),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_15_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(15)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(15),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_14_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(14)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(14),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_14_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(14)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(14),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_13_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(13)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(13),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_13_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(13)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(13),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_12_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(12)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(12),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_12_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(12)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(12),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_11_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(11)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(11),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_11_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(11)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(11),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_10_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(10)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(10),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_10_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(10)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(10),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_9_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(9)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(9),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_9_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(9)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(9),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_8_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(8)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(8),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_8_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(8)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(8),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_7_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(7)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(7),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_7_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(7)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(7),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_6_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(6)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(6),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_6_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(6)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(6),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_5_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(5)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(5),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_5_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(5)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(5),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_4_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(4)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(4),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_4_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(4)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(4),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_3_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(3)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(3),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_3_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(3)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(3),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_2_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(2)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(2),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(2)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(2),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_1_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(1)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(1),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(1),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_0_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => s_axis_divisor_tdata(26),
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(0),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => s_axis_divisor_tdata(26),
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(0),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(26)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(25)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(24)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(23)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(22)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(21)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(20)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(19)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(18)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(17)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(16)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(15)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(14)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(13)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(12)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(11)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(10)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(9)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_q_int(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_27_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_26_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_25_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_24_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_23_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_22_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_21_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_20_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_19_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_18_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_17_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_16_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_15_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_14_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_13_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_12_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_11_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_10_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_9_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_8_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_7_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_6_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_5_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_4_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_3_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_2_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_27_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_26_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_25_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_24_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_23_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_22_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_21_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_20_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_19_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_18_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_17_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_16_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_15_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_14_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_13_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_12_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_11_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_10_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_9_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_8_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_7_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_6_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_5_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_4_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_3_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_2_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(26)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(25)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(24)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(23)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(22)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(21)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(20)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(19)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(18)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(17)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(16)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(15)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(14)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(13)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(12)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(11)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(10)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(9)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_a
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_b
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_int

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_op_a
,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_0_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_0_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_int_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_1_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_1_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_1_MUX_OP_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_2_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_2_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_2_MUX_OP_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_3_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_0_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_0_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_0_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_1_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_1_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_2_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_2_Q
,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP : 
MUXF7
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_3_Q
,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_NO_RTL_USE_MUX7_W_MUX_3_MUX_OP_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_int
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_0_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_int_2_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_OP_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_int_0_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_OP_DEL_RTL_delay_0_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_A_Z_DET_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_all_bits_zero_del
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_A_Z_DET_RTL_delay_0_0_893

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_7_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(7)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_6_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(6)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_5_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(5)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_4_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(4)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_3_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(3)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(2)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => N0,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_7_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_6_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_5_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_4_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_3_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_2_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_1_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_CHAIN_GEN_0_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_1_carry(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_5_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(5)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(13)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_4_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(4)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_3_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(3)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(2)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => N0,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_5_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_4_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_3_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_2_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_1_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_CHAIN_GEN_0_NO_RLOCS_CARRYS_DEL_NEED_DEL_CARRYS_FD : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ZERO_DET_CC_2_CC_carry(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_carry(2)
,
      DI => N0,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_a_ip(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_round_rnd1

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => N0,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX_rt_2543
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_12_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(12)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_12_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(12)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_carry_rnd2

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_11_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(11)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_11_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(11)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_10_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(10)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_10_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(10)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_9_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(9)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_9_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(9)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_8_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(8)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_8_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(8)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_7_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(7)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_7_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(7)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_6_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(6)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_6_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(6)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_5_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(5)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_5_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(5)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_4_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(4)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_4_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(4)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_3_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(3)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_3_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(3)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_2_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(2)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(2)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_1_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(1)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_0_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_round_rnd1
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_round_rnd1
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(12)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(11)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(10)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(9)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_q_int(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_13_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(13)
,
      LI => N0,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_12_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(12)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_12_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(12)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_11_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(11)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_11_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(11)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_10_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(10)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_10_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(10)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_9_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(9)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_9_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(9)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_8_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(8)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_8_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(8)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_7_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(7)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_7_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(7)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_6_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(6)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_6_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(6)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_5_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(5)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_5_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(5)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_4_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(4)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_4_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(4)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_3_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(3)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_3_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(3)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_2_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(2)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_2_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(2)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_1_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(1)
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_1_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(1)
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_0_NO_RLOCS_Q_XOR_SUM_XOR : 
XORCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_carry_rnd2
,
      LI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX : 
MUXCY
    port map (
      CI => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_carry_rnd2
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      S => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_carry(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(13)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(12)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(11)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(10)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(9)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_q_int(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_25 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_25_GND_233_o_MUX_177_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_24 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_24_GND_233_o_MUX_228_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_23 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_23_GND_233_o_MUX_229_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_22 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_22_GND_233_o_MUX_230_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_21 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_21_GND_233_o_MUX_231_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_20 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_20_GND_233_o_MUX_232_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_19 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_19_GND_233_o_MUX_233_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_18 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_18_GND_233_o_MUX_234_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_17 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_17_GND_233_o_MUX_235_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_16 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_16_GND_233_o_MUX_236_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_15 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_15_GND_233_o_MUX_237_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_14 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_14_GND_233_o_MUX_238_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_13 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_13_GND_233_o_MUX_239_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_12 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_12_GND_233_o_MUX_240_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_11 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_11_GND_233_o_MUX_241_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_10 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_10_GND_233_o_MUX_242_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_9 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_9_GND_233_o_MUX_243_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_8 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_8_GND_233_o_MUX_244_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_7 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_7_GND_233_o_MUX_245_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_6 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_6_GND_233_o_MUX_246_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_5 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_5_GND_233_o_MUX_247_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_4 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_4_GND_233_o_MUX_248_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_3 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_3_GND_233_o_MUX_249_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_2 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_2_GND_233_o_MUX_250_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_1 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_1_GND_233_o_MUX_251_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_0 : 
FD
    port map (
      C => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_0_GND_233_o_MUX_252_o
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_div_by_zero_del_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_div_by_zero_del_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout1(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout1(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout2(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout2(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_coarse_est_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_est_prescale_balance_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_use_DSP48E_appDSP48E_0_bppDSP48E_0_need_output_delay_output_delay_dout_i_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_prescaler_gEMBEDDED_MULT_gEMB_MULTS_only_gDSP_iDSP_pi(0, 0, 0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 6),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_0_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_1_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(26),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_28_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_27_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_26_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_25_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_24_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_23_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_22_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_21_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_20_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_19_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_18_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_17_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_16_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_40_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_39_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_38_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_37_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_36_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_35_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_34_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_33_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_32_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_31_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_30_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_29_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_28_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_27_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_26_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_25_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_24_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_23_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_22_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_21_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_20_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_19_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_18_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_17_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_16_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_89 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_89_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_88 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_88_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_88_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_87 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_87_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_87_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_86 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_86_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_86_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_85 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_85_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_85_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_84 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_84_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_84_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_83 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_83_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_83_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_82 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_82_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_82_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_81 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_81_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_81_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_80 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_80_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_80_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_79 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_79_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_79_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_78 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_78_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_78_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_77 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_77_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_77_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_76 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_76_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_76_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_75 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_75_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_75_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_74 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_74_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_74_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_73 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_73_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_73_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_72 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_72_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_72_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_71 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_71_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_71_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_70 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_70_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_70_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_69 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_69_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_69_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_68 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_68_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_68_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_67 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_67_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_67_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_66 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_66_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_66_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_65 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_65_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_65_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_64 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_64_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_64_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_63 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_63_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_63_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_62 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_62_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_62_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_61 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_61_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_61_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_60 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_60_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_60_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_59 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_59_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_59_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_58 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_58_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_58_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_57 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_57_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_57_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_56 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_56_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_56_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_55 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_55_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_55_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_54 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_54_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_54_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_53 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_53_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_53_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_52_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_51 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_51_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_51_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_50 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_50_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_50_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_49 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_49_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_49_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_48 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_48_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_48_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_47 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_47_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_47_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_46 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_46_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_46_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_45 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_45_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_45_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_44 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_44_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_44_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_43 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_43_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_43_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_42 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_42_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_42_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_41 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_41_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_41_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_40 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_40_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_40_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_39 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_39_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_39_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_38 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_38_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_38_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_37_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_37_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_36_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_36_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_35_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_35_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_34_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_34_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_33_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_33_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_32_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_32_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_31_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_31_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_30_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_30_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_29_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_28_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_27_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_26_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_25_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_24_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_23_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_22_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_21_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_20_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_19_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_18_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_17_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_16_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_26 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_27 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(27)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_28 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(28)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_est_reg_opt_has_pipe_first_q_29 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(29)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_subtract_reg_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_subtract_reg_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_subtract_reg_opt_has_pipe_pipe_2_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_subtract_reg_opt_has_pipe_first_q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 14),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 13),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 12),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 11),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 10),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 9),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 8),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 7),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 6),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 14),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 13),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 12),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 11),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 10),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 9),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 8),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 7),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 6),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 14),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 13),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 12),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 11),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 10),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 9),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 8),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 7),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 6),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_14_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_13_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_12_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_11_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_10_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_9_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_8_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_7_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_6_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_5_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_4_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_3_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_2_top_digit_i_extra_digit_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_2_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_pp_digit_i_extra_pp_digit_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_carrysave_del_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_carrysave_del_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_carrysave_del_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denommux_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denommux_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denommux_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_carrysave_carousel_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_47 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_47_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_46 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_46_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_45 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_45_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_44 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_44_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_43 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_43_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_42 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_42_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_41 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_41_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_40 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_40_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_39 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_39_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_38 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_38_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_37_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_36_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_35_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_34_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_33_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_31_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_30_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_29_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_28_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_27_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_26_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_25_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_24_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_23_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_22_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_21_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_20_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_19_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_18_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_17_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_14_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_13_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_12_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_11_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_10_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_9_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_8_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_7_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_6_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_5_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_4_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_3_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_2_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_1_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_residue_reg_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_0_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_32_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_31_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_30_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_29_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_28_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_27_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_26_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_25_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_24_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_23_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_22_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_21_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_20_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_19_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_18_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_17_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_15_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_14_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_13_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_12_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_11_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_10_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_9_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_8_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_7_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_6_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_5_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_4_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_3_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_2_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_1_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_residue_reg_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_0_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_47 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(47)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(47)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_46 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(46)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(46)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_45 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(45)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(45)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_44 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(44)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(44)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_43 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(43)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(43)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_42 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(42)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(42)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_41 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(41)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(41)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_40 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(40)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(40)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_39 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(39)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(39)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_38 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(38)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(38)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(37)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(37)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(36)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(36)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(35)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(35)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(34)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(34)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(33)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(33)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(32)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(32)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(31)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(31)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(30)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(30)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(29)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(29)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(28)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(28)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(27)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(27)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(26)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(25)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(24)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(23)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(22)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(21)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(20)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(19)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(18)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(17)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(16)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(15)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(14)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(13)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(12)
,
      Q => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(11)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(10)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(9)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(8)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(7)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(6)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(5)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(4)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(3)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(2)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(1)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_47 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(47)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_46 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(46)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_45 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(45)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_44 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(44)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_43 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(43)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_42 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(42)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_41 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(41)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_40 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(40)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_39 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(39)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_38 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(38)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(37)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(36)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(35)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(34)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(33)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(32)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(31)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(30)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(29)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(28)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(27)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_digit_balance_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(33)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(33)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(32)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(32)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(31)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(31)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(30)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(30)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(29)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(29)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(28)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(28)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(27)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(27)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(26)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(25)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(24)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(23)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(22)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(21)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(20)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(19)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(18)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(17)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(16)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(15)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(14)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(13)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(12)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(11)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(10)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(9)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(8)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(7)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(6)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(5)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(4)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(3)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(2)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(1)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_quot_carousel_balance_opt_has_pipe_first_q_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(0)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(0)
    );
  U0_i_synth_rdy_if1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_39_135,
      O => m_axis_dout_tvalid
    );
  U0_i_synth_valid_access_in1 : LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_s_axis_dividend_tready,
      I2 => s_axis_dividend_tvalid,
      I3 => s_axis_divisor_tvalid,
      O => U0_i_synth_valid_access_in
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_Mmux_negate_mux11 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(0),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_pipe_4_418
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_pipe_10_688,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT13 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT21 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(11),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT31 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(2),
      I2 => U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT51 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(10),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT61 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(9),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT71 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(8),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT81 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(7),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT91 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(6),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT101 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(5),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT111 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(4),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mmux_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT121 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(3),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line_1_GND_29_o_mux_3_OUT_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm_3_1 : 
LUT4
    generic map(
      INIT => X"5559"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm_4_1 : 
LUT5
    generic map(
      INIT => X"33333363"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm_5_1 : 
LUT5
    generic map(
      INIT => X"FFFFFFFB"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_0_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_18_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_20_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_10_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_12_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_16_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_14_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_16_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_20_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_18_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_2_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_2_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_4_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_8_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_14_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_6_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_8_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_12_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_10_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_1_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_3_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_1_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_11_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_13_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_15_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_17_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_17_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_19_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_19_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_21_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_21_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_3_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_3_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_5_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_5_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_9_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_15_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_7_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_9_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_13_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_7_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_2_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(17)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(9)
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(25)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_3_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(16)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(0)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(8)
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(24)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_1_1 : 
LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(18)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(2)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(10)
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(26)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Madd_EXP_OUT_lut_0_11 : 
LUT3
    generic map(
      INIT => X"41"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Madd_EXP_OUT_lut(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_4_1 : 
LUT5
    generic map(
      INIT => X"44144444"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(4)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(3)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_bdd0
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_5_1 : 
LUT6
    generic map(
      INIT => X"5050505014505050"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(3)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(5)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(2)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(4)
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_bdd0
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_1_1 : 
LUT4
    generic map(
      INIT => X"4414"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(1)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_11 : 
LUT3
    generic map(
      INIT => X"DF"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(1)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_bdd0
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Msub_exp_norm_xor_2_11 : 
LUT3
    generic map(
      INIT => X"59"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_0_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Msub_exp_norm_xor_1_11 : 
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_DIST_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a110 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(0),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a21 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(1),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a31 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(10),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a41 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(11),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a51 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(12),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a61 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(13),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a71 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(14),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a81 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(15),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a91 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(16),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a101 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(17),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a111 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(18),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a121 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(19),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a131 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(2),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a141 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(20),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a151 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(21),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a161 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(22),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a171 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(23),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a181 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(24),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a191 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(25),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a221 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(3),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a231 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(4),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a241 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(5),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a251 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(6),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a261 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(7),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a271 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(8),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Mmux_xor_a281 : 
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(9),
      I1 => s_axis_divisor_tdata(26),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_xor_a(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_a11 : 
LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(19)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_a21 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(25)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(17)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_a31 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(23)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(15)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_a41 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(21)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(13)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_a_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_b11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(11)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_b21 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(9)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_b31 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_Mmux_op_b41 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_op_b_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_a11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_a21 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_1_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_5_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_a31 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_6_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_a41 : 
LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_a_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_b11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_8_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_12_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_b21 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_9_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_13_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_Mmux_op_b31 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_10_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_op_b_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_Mmux_dist_int_1_11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_Mmux_dist_int_3_11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_Mmux_op_a11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_0_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_2_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_a

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_Mmux_op_b11 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_6_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_op_b

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_Mmux_op_a11 : 
LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_Z_op_a

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_all_bits_zero_del1 : 
LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_13_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_all_bits_zero_del

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_1_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(25)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(24)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_2_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(23)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(22)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_3_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(21)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(20)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_4_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(19)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(18)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_5_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(17)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(16)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_6_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(15)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(14)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_7_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(13)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_8_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(11)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_9_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(9)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_10_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(7)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_11_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(5)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_12_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(3)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_13_1 : 
LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(1)
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_a_ip_2_1 : 
LUT3
    generic map(
      INIT => X"7F"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_a_ip(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd214 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_14_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_13_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd221 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_13_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_12_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd231 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_3_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd241 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_2_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd251 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_1_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd261 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_12_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_11_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd271 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_11_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_10_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd281 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_10_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_9_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd291 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_9_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_8_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd2101 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_8_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_7_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd2111 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_7_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_6_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd2121 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_5_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd2131 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_5_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_4_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd2(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1_0_1 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd121 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_26_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_25_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd131 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_17_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_16_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd141 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_16_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_15_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd151 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_15_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_14_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd161 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_25_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_24_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd171 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_24_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_23_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd181 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_23_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_22_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd191 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_22_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_21_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd1101 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_21_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_20_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd1111 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_20_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_19_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd1121 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_19_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_18_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_Mmux_LOGIC_mant_shifted_rnd1131 : 
LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_18_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_17_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_mant_shifted_rnd1(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_0_GND_233_o_MUX_252_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(0)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_0_GND_233_o_MUX_252_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_1_GND_233_o_MUX_251_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(1)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_1_GND_233_o_MUX_251_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_2_GND_233_o_MUX_250_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(2)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_2_GND_233_o_MUX_250_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_4_GND_233_o_MUX_248_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(4)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_4_GND_233_o_MUX_248_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_5_GND_233_o_MUX_247_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(5)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_5_GND_233_o_MUX_247_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_3_GND_233_o_MUX_249_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(3)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_3_GND_233_o_MUX_249_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_6_GND_233_o_MUX_246_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(6)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_6_GND_233_o_MUX_246_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_7_GND_233_o_MUX_245_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(7)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_7_GND_233_o_MUX_245_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_9_GND_233_o_MUX_243_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(9)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_9_GND_233_o_MUX_243_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_10_GND_233_o_MUX_242_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(10)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_10_GND_233_o_MUX_242_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_8_GND_233_o_MUX_244_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(8)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_8_GND_233_o_MUX_244_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_11_GND_233_o_MUX_241_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(11)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_11_GND_233_o_MUX_241_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_12_GND_233_o_MUX_240_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(12)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND1_Q_DEL_RTL_delay_0(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_12_GND_233_o_MUX_240_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_14_GND_233_o_MUX_238_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(14)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_14_GND_233_o_MUX_238_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_15_GND_233_o_MUX_237_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(15)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_15_GND_233_o_MUX_237_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_13_GND_233_o_MUX_239_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(13)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_13_GND_233_o_MUX_239_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_16_GND_233_o_MUX_236_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(16)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_16_GND_233_o_MUX_236_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_17_GND_233_o_MUX_235_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(17)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_17_GND_233_o_MUX_235_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_19_GND_233_o_MUX_233_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(19)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_19_GND_233_o_MUX_233_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_20_GND_233_o_MUX_232_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(20)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_20_GND_233_o_MUX_232_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_18_GND_233_o_MUX_234_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(18)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_18_GND_233_o_MUX_234_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_21_GND_233_o_MUX_231_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(21)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(8)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_21_GND_233_o_MUX_231_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_22_GND_233_o_MUX_230_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(22)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(9)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_22_GND_233_o_MUX_230_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_24_GND_233_o_MUX_228_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(24)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(11)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_24_GND_233_o_MUX_228_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_25_GND_233_o_MUX_177_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(25)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(12)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_25_GND_233_o_MUX_177_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_Mmux_mant_op_23_GND_233_o_MUX_229_o11 : 
LUT4
    generic map(
      INIT => X"4E44"
    )
    port map (
      I0 => aclken,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(23)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(10)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op_23_GND_233_o_MUX_229_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_rfd_i_5_1 : LUT5
    generic map(
      INIT => X"00000001"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_20_Q,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_16_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(8),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(4),
      O => NlwRenamedSig_OI_s_axis_dividend_tready
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_371 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_41_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_381 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_42_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_391 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_43_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_401 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_44_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_411 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_45_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_421 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_46_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_431 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_47_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_331 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_38_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_341 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_39_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_361 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_40_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_321 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_37_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_261 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_251 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_271 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_231 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_611 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_63_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_261 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_601 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_62_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_251 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_591 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_61_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_231 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_581 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_60_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_221 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_561 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_59_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_211 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_551 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_58_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_201 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_541 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_57_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_191 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_181 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_171 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_161 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_151 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_141 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_121 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_111 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_101 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_91 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_711 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_72_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_361 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_40_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_701 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_71_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_341 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_39_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_691 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_70_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_331 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_38_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_671 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_69_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_321 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_37_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_661 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_68_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_311 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_36_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_651 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_67_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_301 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_35_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_641 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_66_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_291 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_34_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_631 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_65_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_281 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_33_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_621 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_64_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_271 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_91 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_141 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_81 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_401 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_71 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_391 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_61 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_421 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_51 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_411 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_8_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_221 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_311 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_28_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_36_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_211 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_301 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_27_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_35_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_201 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_291 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_26_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_34_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_191 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_281 : LUT5
    generic map(
      INIT => X"F7D5A280"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_25_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_33_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_181 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_12_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_171 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_121 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_15_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_161 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_111 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_14_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_101 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_151 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_9_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_13_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_81 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(13),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(15),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(14),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_91 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(14),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(16),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(15),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_71 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(12),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(14),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(13),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_61 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(11),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(13),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(12),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_51 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(10),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(12),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(11),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_41 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(9),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(11),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(10),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_31 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(8),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(10),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(9),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_301 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(7),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(9),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(8),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_291 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(6),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(8),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(7),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_281 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(5),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(7),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(6),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_271 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(4),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(6),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(5),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_261 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(3),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(5),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(4),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_251 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(2),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(4),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(3),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_241 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(1),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(3),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(2),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_131 : LUT5
    generic map(
      INIT => X"E6C4A280"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(2),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(1),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_191 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(23),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(25),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(24),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_211 : LUT5
    generic map(
      INIT => X"FBEA5140"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(25),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(24),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(26),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_201 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(24),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(26),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(25),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_181 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(22),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(24),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(23),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_171 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(21),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(23),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(22),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_151 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(19),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(21),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(20),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_161 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(20),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(22),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(21),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_141 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(18),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(20),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(19),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_121 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(17),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(19),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(18),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_111 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(16),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(18),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(17),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_101 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(15),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(17),
      I4 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(16),
      I5 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_221 : LUT4
    generic map(
      INIT => X"ABA8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(26),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_351 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_4_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_381 : LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_41 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_11_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_7_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_31 : LUT5
    generic map(
      INIT => X"76325410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_10_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_6_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_21 : LUT4
    generic map(
      INIT => X"A820"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(0),
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_11 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_21 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_31 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_41 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_51 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_61 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_71 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_81 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_131 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_241 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_351 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_461 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_571 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_681 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_791 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_901 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_11 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_21 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_131 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_3_41_0_241 : LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_3_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_ctrl_opt_has_pipe_first_q_2_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_2_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_3_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_1_29_0_11 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_1_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_110 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_31 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_41 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_51 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_61 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_71 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_81 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_121 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_171 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_181 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_0_191 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(0, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate11 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(10),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(11),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(12),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(13),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(14),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate91 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_17_1 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(2),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate241 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(3),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate251 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(4),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate261 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(5),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate271 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(6),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate281 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(7),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate291 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(8),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_quot_estimate301 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(9),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux19 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(0),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux21 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(1),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux31 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(10),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux41 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(11),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux51 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(12),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux61 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(13),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux71 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(14),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux81 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(15),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux91 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(16),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux101 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(17),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux111 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(2),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux121 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(3),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux131 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(4),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux141 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(5),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux151 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(6),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux161 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(7),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux171 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(8),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digits_carrysave_mux181 : 
LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(9),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_mux(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_18 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_0_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_37_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_9_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_46_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_10_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_47_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_11_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_48_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_12_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_49_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_13_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_50_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_14_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_51_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom_2_16_1 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_15_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_101 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_1_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_38_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_2_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_39_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_3_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_40_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_4_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_5_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_42_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_151 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_6_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_43_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_161 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_7_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_44_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_2_171 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_8_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_45_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(2, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_17 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_0_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_9_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_30_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_10_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_31_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_11_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_32_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_12_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_33_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_13_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_34_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_14_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_35_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_15_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_36_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_91 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_1_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_101 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_2_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_3_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_4_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_5_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_6_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_27_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_151 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_7_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_28_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_1_161 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_8_Q,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(1, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_17 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_31 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_41 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_51 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_61 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_71 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_81 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_121 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_denom_0_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_denom(0, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_15 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_8_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_9_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_10_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_11_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_12_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_13_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_91 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_101 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_2_141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_7_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_2_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux110 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(10),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(11),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(12),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(13),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(14),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(15),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux91 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(16),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux101 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(17),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(18),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(2),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(3),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(4),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux151 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(5),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux161 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(6),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux171 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(7),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux181 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(8),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_estimate_mux191 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(9),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_mux(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_17 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_31 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_41 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_51 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_61 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_71 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_81 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_121 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_0_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(0, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_17 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_0_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_21 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_1_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_10_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_11_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_12_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_13_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_14_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(26),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_15_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(27),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_91 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_2_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_101 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_3_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_4_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_5_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_6_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_7_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_151 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_8_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_2_161 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_9_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(2, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_17 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_31 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_10_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_41 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_11_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_51 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_12_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_61 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_13_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_71 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_14_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_81 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_15_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_111 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_4_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_121 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_5_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_131 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_6_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_141 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_7_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_151 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_8_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_fb_denom_1_161 : LUT3
    generic map(
      INIT => X"E4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_9_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_scaledenom(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_fb_denom(1, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_110 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_31 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_41 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_51 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_61 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_71 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_81 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_121 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_171 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_181 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_2_191 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(2, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_110 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_21 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_31 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_41 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_51 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_61 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_71 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_81 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_121 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_171 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_181 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_carrysave_1_191 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_carrysave(1, 9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_11 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_21 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_31 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_41 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_51 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_61 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_digit_mux_1_13_0_71 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_mux_1_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_110 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_37_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_27 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_38_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_31 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_47_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_41 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_48_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_51 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_49_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_61 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_50_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_71 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_51_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_131 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_39_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_241 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_40_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_351 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_441 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_42_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_451 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_43_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_461 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_44_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_471 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_45_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_481 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_46_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_110 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_210 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_33 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_31_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_41 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_32_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_51 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_33_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_61 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_34_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_71 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_35_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_81 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_36_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_91 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_101 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_111 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_121 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_131 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_141 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_151 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_161 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_171 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_181 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(26),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_191 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(27),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_201 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(28),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_211 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(29),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_221 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(30),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_231 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_241 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(31),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_251 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(32),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_261 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(33),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_271 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_281 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_291 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_27_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_301 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_28_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_311 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_1_321 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_30_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_1_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_subtract11 : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(18),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_5 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_4 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_3 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_2 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_1 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op_0 : 
FDE
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_Madd_EXP_OUT_lut(0)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX_rt : 
LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_DEL_SHIFT_RTL_delay_0_27_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_RND_BIT_GEN_MODE_NO_NORM_1_OR_0_STRUCT_REQ_GENERAL_LUT6_CHAIN_RND1_CHAIN_GEN_0_NO_RLOCS_C_MUX_CARRY_MUX_rt_2543

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux15 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux21 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_9_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux31 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_10_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux41 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_11_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux51 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_12_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux61 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_13_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux71 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux81 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux91 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux101 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux111 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux121 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux131 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_7_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_i_extra_digits_extra_pp_digit_mux141 : LUT5
    generic map(
      INIT => X"EA404040"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_8_Q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_mux(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_24_1 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp111 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(9)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp91 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(11)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_1_shifted_temp191 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp121 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(8)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp101 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(10)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp51 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(15)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp61 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(14)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp71 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(13)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp81 : 
LUT4
    generic map(
      INIT => X"5410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(12)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_1_shifted_temp201 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_1_shifted_temp211 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp141 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp151 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp161 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp181 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp191 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp171 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp201 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp211 : 
LUT3
    generic map(
      INIT => X"10"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_731 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_74_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_741 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_27_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_75_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_751 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_28_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_76_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_761 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_29_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_77_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_771 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_30_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_78_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_781 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_31_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_79_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_801 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_80_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_811 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_81_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_821 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_82_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_831 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_83_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_841 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_84_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_861 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_86_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_871 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_87_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_851 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_85_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_881 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_88_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_721 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_73_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_22_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_24_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_26_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_23_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_1_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_0_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_25_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_MUX_Z_OP_DEL_RTL_delay_0_2_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_DEL_SHIFT_RTL_delay_0_27_Q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_1_shifted_temp_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_10_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(17)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(9)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(1)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_11_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(16)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(8)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_8_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(19)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(11)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(3)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_9_1 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(18)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(10)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(2)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp231 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(23)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(15)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(7)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp241 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(22)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(14)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(6)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp251 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(21)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(13)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(5)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_Mmux_MUX_LOOP_0_shifted_temp261 : 
LUT6
    generic map(
      INIT => X"5410FEBA54105410"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_3_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(20)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(12)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_c_int_11_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_Z_C_DEL_RTL_delay_0(4)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_NORM_SHIFT_MUX_LOOP_0_shifted_temp_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_531 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_24_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_8_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_40_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_56_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_521 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_23_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_7_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_39_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_55_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_511 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_22_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_6_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_38_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_54_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_501 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_21_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_5_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_37_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_53_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_491 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_20_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_4_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_36_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_52_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_481 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_19_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_3_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_35_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_51_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_471 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_18_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_2_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_34_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_50_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_451 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_17_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_1_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_33_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_49_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_Mmux_shift_mux_5_89_0_441 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_5_Q
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_ctrl_opt_has_pipe_first_q_4_Q
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_16_Q
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_0_Q
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_32_Q
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_4_i_shift_data_opt_has_pipe_first_q_41_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_mux_5_48_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_2_2 : 
LUT5
    generic map(
      INIT => X"44144444"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(2)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(1)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp_3_1 : 
LUT6
    generic map(
      INIT => X"5050505014505050"
    )
    port map (
      I0 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987
,
      I1 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(2)
,
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(3)
,
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(1)
,
      I4 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_EXP_MOD_DEL_RTL_delay_0(0)
,
      I5 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_ROUND_LOGIC_RND2_Q_DEL_RTL_delay_0(13)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_op_exp(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_15_1 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I2 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_101 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_19_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_111 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_20_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_121 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_21_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_141 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_22_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_151 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_23_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_161 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_24_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_171 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_25_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_181 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_26_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_191 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_27_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_201 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_28_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_211 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_29_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_221 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_30_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_231 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_31_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_29_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_251 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_32_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_30_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_Mmux_mux_ab_2_261 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_33_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_31_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_1 : LUT4
    generic map(
      INIT => X"E444"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_47_Q,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate_d(0),
      I3 => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_i_layer_6_i_shift_data_opt_has_pipe_first_q_52_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_mux_ab_2_32_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_BYPASS_INV_403_o1_INV_0 : 
INV
    port map (
      I => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_bypass_balance_opt_has_pipe_first_q
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_BYPASS_INV_403_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_BYPASS_INV_400_o1_INV_0 : 
INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(0),
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_BYPASS_INV_400_o

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_pre_del_offset_16_1_INV_0 : INV
    port map (
      I => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(16)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_pre_del_offset(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero_0_1_INV_0 : 
INV
    port map (
      I => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_M_ABS_Q_DEL_RTL_delay_0(26)
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_chunk_is_zero(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_dist_int_del_4_1_INV_0 : 
INV
    port map (
      I => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_1_MUX_0_OP_DEL_RTL_delay_0_0_1080
,
      O => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_exp_norm(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_0_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_1_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_2_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_3_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_4_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel_0_6_1_5_1_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_prenormalizer_shift_sel(0, 6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim : RAMB16
    generic map(
      DOA_REG => 1,
      DOB_REG => 1,
      INITP_00 => X"AAAAAAAAAAAAAAAAAAAAAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
      INITP_01 => X"5555555555555555555555555555555555555555556AAAAAAAAAAAAAAAAAAAAA",
      INITP_02 => X"0000000000000000000000000000000000000015555555555555555555555555",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"775FD7D777D5FFF77FDFF757D557DD77F77F7FF55F755D5D7F5F75F775D5DD55",
      INITP_05 => X"5F5D5757DDD5DFD577DF5D7D55F75F5F777D55D5DFD7FDFFD775F5FFDDDF5F5F",
      INITP_06 => X"75757DD5D5755DFD7FF7557755777D57F777DF57FD57F5D7775FFD77F7DD75DF",
      INITP_07 => X"7D7D7DD77755F5DFDD77F5F77D55F7F7F55575755FD7555F7DFD5FDFD5FF5575",
      INIT_00 => X"C3D3C799CB64CF32D303D6D9DAB2DE8FE26FE654EA3CEE29F219F60DFA05FE01",
      INIT_01 => X"894E8CDC906E9403979C9B389ED7A27AA621A9CAAD78B129B4DDB895BC51C010",
      INIT_02 => X"5222557D58DB5C3C5FA16308667369E16D5270C6743D77B87B367EB7823B85C3",
      INIT_03 => X"1E072133246227932AC82DFF3139347637B73AF93E3F418844D448234B754ECA",
      INIT_04 => X"ECBEEFBFF2C2F5C8F8D0FBDBFEE901F9050C08220B3A0E561174149417B81ADE",
      INIT_05 => X"BE0EC0E6C3C1C69EC97ECC61CF45D22CD516D802DAF1DDE2E0D6E3CCE6C5E9C0",
      INIT_06 => X"91C39476972C99E49C9E9F5BA21AA4DBA79EAA64AD2CAFF6B2C3B592B864BB37",
      INIT_07 => X"67AF6A406CD46F697201749B773679D47C747F1781BB8461870A89B58C628F11",
      INIT_08 => X"3FA9421B448E4704497B4BF54E7050ED536D55EE58715AF65D7E60076292651F",
      INIT_09 => X"198B1BE01E36208D22E7254227A029FF2C5F2EC23127338D35F5385F3ACB3D39",
      INIT_0A => X"F534F76DF9A7FBE3FE21006102A204E40729096F0BB70E01104C129914E81739",
      INIT_0B => X"D284D4A3D6C4D8E6DB0ADD2FDF56E17FE3A9E5D5E802EA31EC61EE94F0C8F2FD",
      INIT_0C => X"B15FB366B56FB779B984BB91BDA0BFB0C1C2C3D5C5E9C7FFCA17CC30CE4AD066",
      INIT_0D => X"91AB939B958E978199769B6D9D649F5DA158A354A551A750A950AB51AD54AF59",
      INIT_0E => X"7350752C770978E87AC77CA97E8B806F8253843A8621880A89F48BE08DCD8FBB",
      INIT_0F => X"563A580259CB5B965D625F2F60FD62CD649E667068436A176BED6DC46F9C7175",
      INIT_10 => X"3A533C093DC03F78413142EC44A74664482249E04BA14D624F2450E852AC5472",
      INIT_11 => X"1F8B212F22D5247B262327CC29752B202CCC2E79302731D73387353836EB389E",
      INIT_12 => X"05CF076308F80A8F0C260DBE0F5710F1128C142815C6176419031AA41C451DE7",
      INIT_13 => X"ED11EE96F01CF1A2F32AF4B2F63CF7C6F951FADEFC6BFDF9FF89011902AA043C",
      INIT_14 => X"D543D6B9D830D9A8DB21DC9ADE15DF90E10DE28AE408E588E708E889EA0BEB8D",
      INIT_15 => X"BE56BFBEC127C291C3FCC568C6D5C842C9B1CB20CC90CE01CF73D0E5D259D3CD",
      INIT_16 => X"A83EA99AAAF6AC53ADB1AF0FB06FB1CFB330B492B5F4B758B8BCBA21BB87BCEE",
      INIT_17 => X"92F19440959096E1983299849AD79C2B9D7F9ED4A02AA181A2D8A431A58AA6E4",
      INIT_18 => X"7E637FA780EB8230837584BB8602874A889389DC8B268C718DBC8F08905591A3",
      INIT_19 => X"6A8B6BC36CFC6E366F7070AB71E773247461759F76DD781C795C7A9D7BDE7D20",
      INIT_1A => X"575F588D59BB5AEA5C1A5D4B5E7C5FAD60E062136347647B65B066E6681C6953",
      INIT_1B => X"44D645FA471F4844496A4A904BB74CDF4E074F2F5059518352AE53D955055632",
      INIT_1C => X"32EA3404351F363B3757387439913AAF3BCD3CEC3E0C3F2C404D416E429143B3",
      INIT_1D => X"219122A323B424C725DA26ED280229162A2B2B412C582D6F2E862F9E30B731D0",
      INIT_1E => X"10C611CE12D813E114EC15F71702180E191A1A271B351C431D511E611F702080",
      INIT_1F => X"008101810282038404860588068B078F089309970A9C0BA20CA80DAF0EB60FBD",
      INIT_20 => X"03B80378033C030402C8028C0250021401D801980158011C00E000A000600040",
      INIT_21 => X"073406FC06C80694065C062405EC05B405800548050C04D4049C0464042803F0",
      INIT_22 => X"0A680A340A0409D409A00970093C090808D808A40870083C080807D407A0076C",
      INIT_23 => X"0D580D2C0D000CD00CA00C740C480C140BE80BBC0B880B580B280AFC0ACC0A98",
      INIT_24 => X"100C0FE40FB80F900F680F380F0C0EE40EBC0E900E600E340E0C0DE00DB00D84",
      INIT_25 => X"128812641240121811EC11C811A411781150112C110010D810B41088105C1034",
      INIT_26 => X"14D814B81490146C144C1424140013DC13B4139013701348132012FC12D812B0",
      INIT_27 => X"16F816D816B81698167416541634161015EC15CC15AC158415641544151C14F8",
      INIT_28 => X"18F418D818B8189818781858183C181C17FC17DC17BC179C177C175C173C171C",
      INIT_29 => X"1ACC1AAC1A941A781A581A381A1C1A0419E419C419AC198C196C195019301910",
      INIT_2A => X"1C801C681C4C1C301C141BFC1BE41BC41BA81B901B741B581B3C1B201B001AE8",
      INIT_2B => X"1E181E001DE81DD01DB81D9C1D841D6C1D501D381D201D041CE81CCC1CB81C9C",
      INIT_2C => X"1F981F801F681F541F3C1F241F081EF01EDC1EC41EAC1E941E7C1E641E4C1E34",
      INIT_2D => X"20FC20E820D020BC20A42090207C2064204C20342020200C1FF41FDC1FC41FAC",
      INIT_2E => X"224C22382220221021F821E421D021BC21A82190217C21682154213C21282110",
      INIT_2F => X"23842374235C234C233C2324231022FC22E822D822C422B0229C22882274225C",
      INIT_30 => X"24A8249C24882474246424502440242C241C240823F423E423D023C023AC2394",
      INIT_31 => X"25C025B025A02590257C256C255C2548253825282514250424F424E024D024BC",
      INIT_32 => X"26C826B826A4269426882678266426542648263426242614260025F425E425D0",
      INIT_33 => X"27B827AC27A0279027802770276027542744273027242714270426F826E426D4",
      INIT_34 => X"28A4289828882878286C286028502840283028242814280427F827E827DC27CC",
      INIT_35 => X"297C2974296829582948293C293029202914290828F828E828DC28D028C028B0",
      INIT_36 => X"2A502A442A382A282A1C2A102A0429F829E829DC29D029C029B429A8299C298C",
      INIT_37 => X"2B142B082AFC2AF02AE42AD82ACC2AC02AB42AA42A9C2A902A802A742A682A5C",
      INIT_38 => X"2BCC2BC42BB82BAC2BA42B982B882B7C2B742B682B582B502B442B382B2C2B20",
      INIT_39 => X"2C802C742C6C2C602C542C482C3C2C342C282C1C2C142C082BFC2BF02BE42BD8",
      INIT_3A => X"2D282D1C2D142D082CFC2CF42CEC2CE02CD42CC82CC02CB82CA82C9C2C942C8C",
      INIT_3B => X"2DC82DBC2DB42DA82DA02D982D882D802D7C2D702D642D582D4C2D482D3C2D30",
      INIT_3C => X"2E602E542E4C2E442E382E302E282E1C2E142E0C2E002DF42DF02DE42DD82DD4",
      INIT_3D => X"2EEC2EE82EE02ED42ECC2EC02EB82EB42EA82E9C2E942E8C2E842E7C2E702E68",
      INIT_3E => X"2F782F702F682F602F542F502F482F3C2F342F2C2F242F1C2F102F082F042EF8",
      INIT_3F => X"2FF82FF42FEC2FE42FDC2FD42FCC2FC42FBC2FB42FAC2FA02F982F942F8C2F80",
      INIT_A => X"000000000",
      INIT_B => X"000000000",
      INIT_FILE => "NONE",
      INVERT_CLK_DOA_REG => FALSE,
      INVERT_CLK_DOB_REG => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      SIM_COLLISION_CHECK => "NONE",
      SRVAL_A => X"000000000",
      SRVAL_B => X"000000000",
      WRITE_MODE_A => "READ_FIRST",
      WRITE_MODE_B => "READ_FIRST",
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 18
    )
    port map (
      CASCADEINA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CASCADEINB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CLKA => aclk,
      CLKB => aclk,
      ENA => aclken,
      REGCEA => aclken,
      REGCEB => aclken,
      ENB => aclken,
      SSRA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      SSRB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CASCADEOUTA => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_CASCADEOUTA_UNCONNECTED
,
      CASCADEOUTB => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_CASCADEOUTB_UNCONNECTED
,
      ADDRA(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRA(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRA(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(25)
,
      ADDRA(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(24)
,
      ADDRA(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(23)
,
      ADDRA(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(22)
,
      ADDRA(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(21)
,
      ADDRA(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(20)
,
      ADDRA(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(19)
,
      ADDRA(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(18)
,
      ADDRA(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(17)
,
      ADDRA(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRA(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRA(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRA(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRB(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRB(13) => N0,
      ADDRB(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(25)
,
      ADDRB(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(24)
,
      ADDRB(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(23)
,
      ADDRB(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(22)
,
      ADDRB(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(21)
,
      ADDRB(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(20)
,
      ADDRB(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(19)
,
      ADDRB(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(18)
,
      ADDRB(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(17)
,
      ADDRB(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRB(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRB(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ADDRB(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIA(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIB(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPA(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPA(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPA(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPA(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPB(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPB(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPB(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DIPB(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEA(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEA(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEA(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEA(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEB(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEB(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEB(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      WEB(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      DOA(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_31_UNCONNECTED
,
      DOA(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_30_UNCONNECTED
,
      DOA(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_29_UNCONNECTED
,
      DOA(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_28_UNCONNECTED
,
      DOA(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_27_UNCONNECTED
,
      DOA(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_26_UNCONNECTED
,
      DOA(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_25_UNCONNECTED
,
      DOA(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_24_UNCONNECTED
,
      DOA(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_23_UNCONNECTED
,
      DOA(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_22_UNCONNECTED
,
      DOA(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_21_UNCONNECTED
,
      DOA(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_20_UNCONNECTED
,
      DOA(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_19_UNCONNECTED
,
      DOA(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_18_UNCONNECTED
,
      DOA(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_17_UNCONNECTED
,
      DOA(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOA_16_UNCONNECTED
,
      DOA(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(15),
      DOA(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(14),
      DOA(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(13),
      DOA(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(12),
      DOA(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(11),
      DOA(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(10),
      DOA(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(9),
      DOA(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(8),
      DOA(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(7),
      DOA(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(6),
      DOA(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(5),
      DOA(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(4),
      DOA(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(3),
      DOA(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(2),
      DOA(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(1),
      DOA(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout1(0),
      DOB(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_31_UNCONNECTED
,
      DOB(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_30_UNCONNECTED
,
      DOB(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_29_UNCONNECTED
,
      DOB(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_28_UNCONNECTED
,
      DOB(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_27_UNCONNECTED
,
      DOB(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_26_UNCONNECTED
,
      DOB(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_25_UNCONNECTED
,
      DOB(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_24_UNCONNECTED
,
      DOB(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_23_UNCONNECTED
,
      DOB(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_22_UNCONNECTED
,
      DOB(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_21_UNCONNECTED
,
      DOB(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_20_UNCONNECTED
,
      DOB(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_19_UNCONNECTED
,
      DOB(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_18_UNCONNECTED
,
      DOB(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_17_UNCONNECTED
,
      DOB(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOB_16_UNCONNECTED
,
      DOB(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(15),
      DOB(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(14),
      DOB(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(13),
      DOB(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(12),
      DOB(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(11),
      DOB(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(10),
      DOB(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(9),
      DOB(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(8),
      DOB(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(7),
      DOB(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(6),
      DOB(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(5),
      DOB(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(4),
      DOB(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(3),
      DOB(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(2),
      DOB(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(1),
      DOB(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(0),
      DOPA(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPA_3_UNCONNECTED
,
      DOPA(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPA_2_UNCONNECTED
,
      DOPA(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout1(1),
      DOPA(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout1(0),
      DOPB(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPB_3_UNCONNECTED
,
      DOPB(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_i_not_sandia_i_prim_DOPB_2_UNCONNECTED
,
      DOPB(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout2(1),
      DOPB(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_parout2(0)
    );
  U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q,
      CE => aclken,
      Q => NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0_Q_UNCONNECTED,
      Q31 => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0_2544,
      A(4) => N0,
      A(3) => N0,
      A(2) => N0,
      A(1) => N0,
      A(0) => N0
    );
  U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_0_2544,
      CE => aclken,
      Q => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1_2545,
      Q31 => NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1_Q31_UNCONNECTED,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(2) => N0,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_39_1_2545,
      Q => U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_39_135
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_first_q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4_2546
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_pipe_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_Mshreg_opt_has_pipe_pipe_4_2546
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_negate_carousel_opt_has_pipe_pipe_4_418

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(26),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26_2547,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_26 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_26_2547,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(25),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25_2548,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_25_2548,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(22),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22_2549,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_22_2549,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(24),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24_2550,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_24_2550,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(23),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23_2551,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_23_2551,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(19),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19_2552,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_19_2552,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(21),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21_2553,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_21_2553,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(20),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20_2554,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_20_2554,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16_2555,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_16_2555,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18_2556,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_18_2556,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17_2557,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_17_2557,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15_2558,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_15_2558,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14_2559,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_14_2559,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13_2560,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_13_2560,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12_2561,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_12_2561,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9_2562,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_9_2562,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11_2563,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_11_2563,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10_2564,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_10_2564,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6_2565,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_6_2565,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8_2566,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_8_2566,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7_2567,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_7_2567,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3_2568,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_3_2568,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5_2569,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_5_2569,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4_2570,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_4_2570,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2_2571,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_2_2571,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1_2572,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_1_2572,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_dividend_tdata(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0_2573,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_Mshreg_opt_has_pipe_pipe_9_0_2573,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_numer_del_opt_has_pipe_pipe_9(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_A_Z_DET_RTL_delay_0_0_893
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1_2574
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_Mshreg_RTL_delay_1_2574
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_EXP_ZERO_DELAY_RTL_delay_1_987

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_16_Q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20_2575,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_20_2575,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_4_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0_2576
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_0_2576
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_norm_dist_skew_3_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1_2577
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_Mshreg_RTL_delay_1_1_2577
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_LZE_ENCODE_0_DIST_DEL_RTL_delay_1_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => s_axis_divisor_tdata(26),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q_2578,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_first_q : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_first_q_2578,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_first_q_1227
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_NEW_CODE_ND_DEL_DEL_GT_1_delay_line(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15_2579,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_Mshreg_nd_pipe_15_2579,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_flow_ctrl_nd_pipe_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(14)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14_2580,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_14_2580,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_pre_del_offset(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16_2581,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_16_2581,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(15)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15_2582,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_15_2582,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(13)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13_2583,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_13_2583,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(12)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12_2584,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_12_2584,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(11)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11_2585,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_11_2585,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(10)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10_2586,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_10_2586,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(7)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7_2587,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_7_2587,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(9)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9_2588,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_9_2588,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(8)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8_2589,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_8_2589,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(4)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4_2590,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_4_2590,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(6)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6_2591,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_6_2591,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(5)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5_2592,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_5_2592,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(1)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1_2593,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_1_2593,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(3)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3_2594,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_3_2594,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(2)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2_2595,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_2_2595,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(0)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0_2596,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_Mshreg_del_addr_offset_0_2596,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => N0,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26_2597,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_26 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_26_2597,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(25)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25_2598,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_25_2598,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(24)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24_2599,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_24_2599,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(21)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21_2600,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_21_2600,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(23)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23_2601,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_23_2601,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(22)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22_2602,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_22_2602,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(18)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18_2603,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_18_2603,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(20)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20_2604,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_20_2604,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(19)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19_2605,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_19_2605,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(17)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17_2606,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_17_2606,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_mant_op(16)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16_2607,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_16_2607,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5_2608,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_5_2608,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4_2609,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_4_2609,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1_2610,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_1_2610,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3_2611,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_3_2611,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2_2612,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_2_2612,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_bypass_balance_opt_has_pipe_first_q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1_2613,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_1_2613,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_fix_to_flt_i_fpo_FLT_PT_OP_FIX_TO_FLT_OP_SPD_OP_OP_exp_op(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0_2614,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_Mshreg_opt_has_pipe_pipe_3_0_2614,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fix_prenorm_i_shift_del_opt_has_pipe_pipe_3(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_first_q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3_2615,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_Mshreg_opt_has_pipe_pipe_3_2615,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_del_opt_has_pipe_pipe_3_2306
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_12_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12_2616
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_12_2616
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_13_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13_2617
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_13_2617
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_9_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9_2618
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_9_2618
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_11_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11_2619
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_11_2619
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_10_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10_2620
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_10_2620
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6_2621
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_6_2621
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_8_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8_2622
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_8_2622
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_first_q_7_Q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7_2623
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_Mshreg_opt_has_pipe_pipe_4_7_2623
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digits_1_lower_digits_i_extra_digit_carousel_opt_has_pipe_pipe_4_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(16),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16_2624
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_16_2624
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18_2625
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_18_2625
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(17),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17_2626
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_17_2626
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(15),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15_2627
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_15_2627
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(14),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14_2628
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_14_2628
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(13),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13_2629
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_13_2629
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(12),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12_2630
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_12_2630
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(9),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9_2631
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_9_2631
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(11),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11_2632
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_11_2632
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(10),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10_2633
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_10_2633
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(6),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6_2634
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_6_2634
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(8),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8_2635
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_8_2635
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(7),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7_2636
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_7_2636
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3_2637
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_3_2637
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(5),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5_2638
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_5_2638
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(4),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4_2639
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_4_2639
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2_2640
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_2_2640
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1_2641
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_1_2641
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_reg_opt_has_pipe_first_q(0),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0_2642
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_Mshreg_opt_has_pipe_pipe_3_0_2642
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_est_carousel_opt_has_pipe_pipe_3(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2643
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2643
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2644
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2644
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2645
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2645
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2646
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2646
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2647
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2647
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2648
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2648
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2649
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2649
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2650
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2650
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2651
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2651
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2652
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2652
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2653
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2653
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2654
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2654
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2655
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2655
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2656
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2656
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2657
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2657
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2658
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2658
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_reg_opt_has_pipe_first_q_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2659
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2659
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_denom_pipe_opt_has_pipe_pipe_3_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2660
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2660
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2661
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2661
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2662
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2662
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2663
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2663
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2664
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2664
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2665
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2665
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2666
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2666
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2667
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2667
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2668
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2668
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2669
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2669
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2670
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2670
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2671
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2671
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2672
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2672
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2673
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2673
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_reg_opt_has_pipe_first_q_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2674
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2674
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_denom_pipe_opt_has_pipe_pipe_3_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_13_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2675
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_13_2675
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_15_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2676
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_15_2676
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_14_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2677
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_14_2677
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_12_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2678
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_12_2678
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_11_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2679
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_11_2679
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_10_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2680
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_10_2680
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_9_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2681
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_9_2681
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_6_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2682
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_6_2682
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_8_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2683
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_8_2683
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_7_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2684
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_7_2684
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_3_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2685
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_3_2685
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_5_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2686
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_5_2686
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_4_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2687
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_4_2687
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_0_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2688
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_0_2688
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_2_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2689
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_2_2689
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_reg_opt_has_pipe_first_q_1_Q,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2690
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_Mshreg_opt_has_pipe_pipe_3_1_2690
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_denom_pipe_opt_has_pipe_pipe_3_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(59),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37_2691
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_37 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_37_2691
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(58),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36_2692
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_36 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_36_2692
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(36)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(57),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35_2693
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_35 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_35_2693
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(35)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(56),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34_2694
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_34 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_34_2694
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(34)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(53),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31_2695
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_31 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_31_2695
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(31)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(55),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33_2696
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_33 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_33_2696
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(33)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(54),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32_2697
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_32 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_32_2697
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(32)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(50),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28_2698
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_28 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_28_2698
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(28)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(52),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30_2699
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_30 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_30_2699
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(30)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(51),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29_2700
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_29 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_29_2700
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(29)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(47),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25_2701
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_25 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_25_2701
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(25)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(49),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27_2702
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_27 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_27_2702
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(27)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(48),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26_2703
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_26 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_26_2703
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(26)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(46),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24_2704
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_24 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_24_2704
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(24)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(45),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23_2705
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_23 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_23_2705
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(23)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(44),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22_2706
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_22 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_22_2706
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(22)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(43),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21_2707
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_21 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_21_2707
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(21)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(40),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18_2708
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_18 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_18_2708
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(18)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(42),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20_2709
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_20 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_20_2709
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(20)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(41),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19_2710
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_19 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_19_2710
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(19)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(37),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15_2711
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_15 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_15_2711
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(15)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(39),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17_2712
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_17 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_17_2712
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(17)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(38),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16_2713
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_16 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_16_2713
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(16)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(46)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12_2714
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_12 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_12_2714
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(12)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => NlwRenamedSig_OI_m_axis_dout_tdata(36),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14_2715
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_14 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_14_2715
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(14)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(47)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13_2716
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_13 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_13_2716
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(13)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(43)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9_2717
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_9 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_9_2717
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(9)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(45)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11_2718
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_11 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_11_2718
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(11)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(44)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10_2719
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_10 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_10_2719
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(10)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(40)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6_2720
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_6 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_6_2720
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(6)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(42)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8_2721
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_8 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_8_2721
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(8)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(41)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7_2722
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_7 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_7_2722
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(7)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(37)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3_2723
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_3 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_3_2723
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(3)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(39)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5_2724
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_5 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_5_2724
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(5)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(38)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4_2725
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_4 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_4_2725
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(4)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(34)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0_2726
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_0 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_0_2726
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(0)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(36)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2_2727
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_2 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_2_2727
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(2)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1 : 
SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => 
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_p_balance_opt_has_pipe_first_q(35)
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1_2728
,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d_1 : 
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_Mshreg_i_vx5_sp3_i_casc_dsp48_OP_A_d_1_2728
,
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(1)

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => N0,
      A2 => N0,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_first_q_1227,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10_2729,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_pipe_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_Mshreg_opt_has_pipe_pipe_10_2729,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_fixed_i_negate_del_opt_has_pipe_pipe_10_688
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15_2730,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_15_2730,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14_2731,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_14_2731,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13_2732,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_13_2732,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12_2733,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_12_2733,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11_2734,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_11_2734,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8_2735,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_8_2735,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10_2736,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_10_2736,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9_2737,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_9_2737,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5_2738,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_5_2738,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7_2739,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_7_2739,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6_2740,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_6_2740,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2_2741,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_2_2741,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4_2742,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_4_2742,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3_2743,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_3_2743,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1_2744,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_1_2744,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => N0,
      A1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0_2745,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_fulldenom_d_0_2745,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_fulldenom_d(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(1),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2_2746,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_2_2746,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(2),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3_2747,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_3_2747,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(3),
      Q => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4_2748,
      Q15 => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4_Q15_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_Mshreg_opt_has_pipe_first_q_4_2748,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A1 => N0,
      A2 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A3 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CE => aclken,
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_nd_pipe2_opt_has_pipe_first_q(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit_2749,
      Q15 => NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit_Q15_UNCONNECTED
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_last_digit : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_Mshreg_last_digit_2749,
      Q => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_last_digit_518
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CLK => aclk,
      CARRYCASCIN => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_carrycascout
,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => N0,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_BYPASS_INV_403_o
,
      OPMODE(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_BYPASS_INV_403_o
,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_negate_balance_opt_has_pipe_first_q
,
      ALUMODE(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_negate_balance_opt_has_pipe_first_q
,
      C(47) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(46) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(45) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(44) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(43) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(42) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(41) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(40) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(39) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(38) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(37) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(37)
,
      C(36) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(36)
,
      C(35) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(35)
,
      C(34) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(34)
,
      C(33) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(33)
,
      C(32) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(32)
,
      C(31) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(31)
,
      C(30) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(30)
,
      C(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(29)
,
      C(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(28)
,
      C(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(27)
,
      C(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(26)
,
      C(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(25)
,
      C(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(24)
,
      C(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(23)
,
      C(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(22)
,
      C(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(21)
,
      C(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(20)
,
      C(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(19)
,
      C(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(18)
,
      C(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(17)
,
      C(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(16)
,
      C(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(15)
,
      C(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(14)
,
      C(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(13)
,
      C(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(12)
,
      C(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(11)
,
      C(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(10)
,
      C(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(9)
,
      C(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(8)
,
      C(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(7)
,
      C(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(6)
,
      C(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(5)
,
      C(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(4)
,
      C(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(3)
,
      C(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(2)
,
      C(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(1)
,
      C(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_OP_A_d(0)
,
      B(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(17)
,
      B(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(16)
,
      B(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(15)
,
      B(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(14)
,
      B(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(13)
,
      B(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(12)
,
      B(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(11)
,
      B(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(10)
,
      B(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(9)
,
      B(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(8)
,
      B(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(7)
,
      B(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(6)
,
      B(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(5)
,
      B(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(4)
,
      B(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(3)
,
      B(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(2)
,
      B(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(1)
,
      B(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(0)
,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => NlwRenamedSignal_m_axis_dout_tdata(72),
      P(35) => m_axis_dout_tdata(71),
      P(34) => m_axis_dout_tdata(70),
      P(33) => m_axis_dout_tdata(69),
      P(32) => m_axis_dout_tdata(68),
      P(31) => m_axis_dout_tdata(67),
      P(30) => m_axis_dout_tdata(66),
      P(29) => m_axis_dout_tdata(65),
      P(28) => m_axis_dout_tdata(64),
      P(27) => m_axis_dout_tdata(63),
      P(26) => m_axis_dout_tdata(62),
      P(25) => m_axis_dout_tdata(61),
      P(24) => m_axis_dout_tdata(60),
      P(23) => NlwRenamedSig_OI_m_axis_dout_tdata(59),
      P(22) => NlwRenamedSig_OI_m_axis_dout_tdata(58),
      P(21) => NlwRenamedSig_OI_m_axis_dout_tdata(57),
      P(20) => NlwRenamedSig_OI_m_axis_dout_tdata(56),
      P(19) => NlwRenamedSig_OI_m_axis_dout_tdata(55),
      P(18) => NlwRenamedSig_OI_m_axis_dout_tdata(54),
      P(17) => NlwRenamedSig_OI_m_axis_dout_tdata(53),
      P(16) => NlwRenamedSig_OI_m_axis_dout_tdata(52),
      P(15) => NlwRenamedSig_OI_m_axis_dout_tdata(51),
      P(14) => NlwRenamedSig_OI_m_axis_dout_tdata(50),
      P(13) => NlwRenamedSig_OI_m_axis_dout_tdata(49),
      P(12) => NlwRenamedSig_OI_m_axis_dout_tdata(48),
      P(11) => NlwRenamedSig_OI_m_axis_dout_tdata(47),
      P(10) => NlwRenamedSig_OI_m_axis_dout_tdata(46),
      P(9) => NlwRenamedSig_OI_m_axis_dout_tdata(45),
      P(8) => NlwRenamedSig_OI_m_axis_dout_tdata(44),
      P(7) => NlwRenamedSig_OI_m_axis_dout_tdata(43),
      P(6) => NlwRenamedSig_OI_m_axis_dout_tdata(42),
      P(5) => NlwRenamedSig_OI_m_axis_dout_tdata(41),
      P(4) => NlwRenamedSig_OI_m_axis_dout_tdata(40),
      P(3) => NlwRenamedSig_OI_m_axis_dout_tdata(39),
      P(2) => NlwRenamedSig_OI_m_axis_dout_tdata(38),
      P(1) => NlwRenamedSig_OI_m_axis_dout_tdata(37),
      P(0) => NlwRenamedSig_OI_m_axis_dout_tdata(36),
      A(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(47)
,
      A(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(46)
,
      A(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(45)
,
      A(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(44)
,
      A(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(43)
,
      A(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(42)
,
      A(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(41)
,
      A(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(40)
,
      A(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(39)
,
      A(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(38)
,
      A(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(37)
,
      A(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(36)
,
      A(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(35)
,
      A(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(34)
,
      A(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(33)
,
      A(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(32)
,
      A(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(31)
,
      A(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(30)
,
      A(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(29)
,
      A(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(28)
,
      A(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(27)
,
      A(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(26)
,
      A(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(25)
,
      A(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(24)
,
      A(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(23)
,
      A(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(22)
,
      A(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(21)
,
      A(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(20)
,
      A(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(19)
,
      A(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_abport2(18)
,
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_upper_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CARRYCASCOUT => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_carrycascout
,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_BYPASS_INV_400_o
,
      OPMODE(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_BYPASS_INV_400_o
,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_negate_mux,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(33),
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(32),
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(31),
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(30),
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(29),
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(28),
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(27),
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(26),
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(25),
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(24),
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(23),
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(22),
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(21),
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(20),
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(19),
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(18),
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(17),
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(16),
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(15),
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(14),
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(13),
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(12),
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(11),
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(10),
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(9),
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(8),
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(7),
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(6),
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(5),
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(4),
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(3),
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(2),
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(1),
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_result_fb(0),
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_last_digit_518,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(14),
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(13),
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(12),
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(11),
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(10),
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(9),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(8),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(7),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(6),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(5),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(4),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(3),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(2),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(1),
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(0),
      P(47) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(47)
,
      P(46) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(46)
,
      P(45) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(45)
,
      P(44) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(44)
,
      P(43) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(43)
,
      P(42) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(42)
,
      P(41) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(41)
,
      P(40) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(40)
,
      P(39) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(39)
,
      P(38) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(38)
,
      P(37) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(37)
,
      P(36) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(36)
,
      P(35) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(35)
,
      P(34) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(34)
,
      P(33) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(33)
,
      P(32) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(32)
,
      P(31) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(31)
,
      P(30) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(30)
,
      P(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(29)
,
      P(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(28)
,
      P(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(27)
,
      P(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(26)
,
      P(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(25)
,
      P(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(24)
,
      P(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(23)
,
      P(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(22)
,
      P(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(21)
,
      P(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(20)
,
      P(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(19)
,
      P(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(18)
,
      P(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(17)
,
      P(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(16)
,
      P(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(15)
,
      P(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(14)
,
      P(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(13)
,
      P(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(12)
,
      P(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(11)
,
      P(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(10)
,
      P(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(9)
,
      P(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(8)
,
      P(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(7)
,
      P(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(6)
,
      P(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(5)
,
      P(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(4)
,
      P(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(3)
,
      P(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(2)
,
      P(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(1)
,
      P(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_pport1(0)
,
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_quotient_collector_i_typical_case_i_addsub_i_vx5_sp3_i_casc_dsp48_i_lower_addsub_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(29) => N0,
      A(28) => N0,
      A(27) => N0,
      A(26) => N0,
      A(25) => N0,
      A(24) => N0,
      A(23) => N0,
      A(22) => N0,
      A(21) => N0,
      A(20) => N0,
      A(19) => N0,
      A(18) => N0,
      A(17) => N0,
      A(16) => N0,
      A(15) => N0,
      A(14) => N0,
      A(13) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(13),
      A(12) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(12),
      A(11) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(11),
      A(10) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(10),
      A(9) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(9),
      A(8) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(8),
      A(7) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(7),
      A(6) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(6),
      A(5) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(5),
      A(4) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(4),
      A(3) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(3),
      A(2) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(2),
      A(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(1),
      A(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_lut_i_synth_opt_i_synth_fullprim_dataout2(0),
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => N0,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(21),
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(20),
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(19),
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(18),
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(17),
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(16),
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(15),
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(14),
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(13),
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(12),
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(11),
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(10),
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(9),
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(8),
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(7),
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(6),
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(5),
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(4),
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(3),
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(2),
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(1),
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_coarse_est_d(0),
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(16),
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(16),
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(15),
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(14),
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(13),
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(12),
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(11),
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(10),
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(9),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(8),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(7),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(6),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(5),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(4),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(3),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(2),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(1),
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_del_addr_offset(0),
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(18),
      P(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(17),
      P(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(16),
      P(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(15),
      P(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(14),
      P(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(13),
      P(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(12),
      P(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(11),
      P(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(10),
      P(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(9),
      P(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(8),
      P(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(7),
      P(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(6),
      P(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(5),
      P(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(4),
      P(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(3),
      P(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(2),
      P(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(1),
      P(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_estimate(0),
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED
,
      P(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED
,
      P(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED
,
      P(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED
,
      P(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED
,
      P(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED
,
      P(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED
,
      P(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED
,
      P(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED
,
      P(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED
,
      P(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED
,
      P(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED
,
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_estimator_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 47),
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 46),
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 45),
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 44),
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 43),
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 42),
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 41),
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 40),
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 39),
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 38),
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 37),
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 36),
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 35),
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 34),
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 33),
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 32),
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 31),
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 30),
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 29),
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 28),
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 27),
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 26),
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 25),
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 24),
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 23),
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 22),
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 21),
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 20),
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 19),
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 18),
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 17),
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 16),
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 15),
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 14),
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 13),
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 12),
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 11),
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 10),
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 9),
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 8),
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 7),
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 6),
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 5),
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 4),
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 3),
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 2),
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 1),
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 0),
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_17_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_16_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_15_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_14_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_13_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_12_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_11_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_10_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_9_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_8_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_7_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_6_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_5_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_4_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_3_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_2_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_2_1_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(15),
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(14),
      P(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(13),
      P(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(12),
      P(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(11),
      P(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(10),
      P(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(9),
      P(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(8),
      P(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(7),
      P(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(6),
      P(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(5),
      P(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(4),
      P(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(3),
      P(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(2),
      P(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(1),
      P(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_quot_digit(0),
      P(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_18_Q,
      P(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_17_Q,
      P(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_16_Q,
      P(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_15_Q,
      P(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_14_Q,
      P(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_13_Q,
      P(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_12_Q,
      P(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_11_Q,
      P(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_10_Q,
      P(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_9_Q,
      P(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_8_Q,
      P(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_7_Q,
      P(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_6_Q,
      P(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_5_Q,
      P(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_4_Q,
      P(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_3_Q,
      P(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_2_Q,
      P(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_1_Q,
      P(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_2_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(29),
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(28),
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(27),
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(26),
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(25),
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(24),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(23),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(22),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(21),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(20),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(19),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(18),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(17),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(16),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(15),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(14),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(13),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(12),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(11),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(10),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(9),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(8),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(7),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(6),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(5),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(4),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(3),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(2),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(1),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 47),
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 46),
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 45),
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 44),
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 43),
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 42),
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 41),
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 40),
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 39),
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 38),
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 37),
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 36),
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 35),
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 34),
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 33),
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 32),
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 31),
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 30),
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 29),
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 28),
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 27),
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 26),
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 25),
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 24),
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 23),
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 22),
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 21),
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 20),
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 19),
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 18),
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 17),
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 16),
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 15),
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 14),
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 13),
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 12),
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 11),
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 10),
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 9),
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 8),
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 7),
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 6),
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 5),
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 4),
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 3),
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 2),
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 1),
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 0),
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_16_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_15_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_14_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_13_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_12_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_11_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_10_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_9_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_8_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_7_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_6_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_5_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_4_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_3_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_2_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_1_1_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_47_Q,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_33_Q,
      P(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_32_Q,
      P(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_31_Q,
      P(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_30_Q,
      P(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_29_Q,
      P(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_28_Q,
      P(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_27_Q,
      P(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_26_Q,
      P(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_25_Q,
      P(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_24_Q,
      P(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_23_Q,
      P(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_22_Q,
      P(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_21_Q,
      P(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_20_Q,
      P(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_19_Q,
      P(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_18_Q,
      P(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_17_Q,
      P(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_16_Q,
      P(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_15_Q,
      P(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_14_Q,
      P(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_13_Q,
      P(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_12_Q,
      P(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_11_Q,
      P(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_10_Q,
      P(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_9_Q,
      P(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_8_Q,
      P(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_7_Q,
      P(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_6_Q,
      P(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_5_Q,
      P(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_4_Q,
      P(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_3_Q,
      P(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_2_Q,
      P(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_1_Q,
      P(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_1_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(29),
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(28),
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(27),
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(26),
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(25),
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(24),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(23),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(22),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(21),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(20),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(19),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(18),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(17),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(16),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(15),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(14),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(13),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(12),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(11),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(10),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(9),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(8),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(7),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(6),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(5),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(4),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(3),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(2),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(1),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 47),
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 46),
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 45),
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 44),
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 43),
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 42),
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 41),
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 40),
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 39),
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 38),
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 37),
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 36),
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 35),
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 34),
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 33),
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 32),
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 31),
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 30),
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 29),
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 28),
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 27),
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 26),
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 25),
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 24),
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 23),
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 22),
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 21),
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 20),
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 19),
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 18),
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 17),
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 16),
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 15),
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 14),
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 13),
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 12),
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 11),
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 10),
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 9),
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 8),
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 7),
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 6),
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 5),
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 4),
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 3),
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 2),
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 1),
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 0),
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_subtract_d,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_16_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_15_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_14_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_13_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_12_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_11_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_10_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_9_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_8_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_7_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_6_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_5_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_4_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_3_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_2_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_denom_d_0_1_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_18_Q,
      P(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_17_Q,
      P(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_16_Q,
      P(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_15_Q,
      P(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_14_Q,
      P(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_13_Q,
      P(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_12_Q,
      P(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_11_Q,
      P(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_10_Q,
      P(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_9_Q,
      P(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_8_Q,
      P(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_7_Q,
      P(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_6_Q,
      P(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_5_Q,
      P(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_4_Q,
      P(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_3_Q,
      P(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_2_Q,
      P(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_1_Q,
      P(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_out_0_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(29),
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(28),
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(27),
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(26),
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(25),
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(24),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(23),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(22),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(21),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(20),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(19),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(18),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(17),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(16),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(15),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(14),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(13),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(12),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(11),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(10),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(9),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(8),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(7),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(6),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(5),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(4),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(3),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(2),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(1),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_quot_estimate_d(0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_mult_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CECTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => N0,
      OPMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(0) => N0,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(47),
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(46),
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(45),
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(44),
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(43),
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(42),
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(41),
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(40),
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(39),
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(38),
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(37),
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(36),
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(35),
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(34),
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(33),
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(32),
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(31),
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(30),
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(29),
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(28),
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(27),
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(26),
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(25),
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(24),
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(23),
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(22),
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(21),
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(20),
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(19),
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(18),
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(17),
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(16),
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(15),
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(14),
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(13),
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(12),
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(11),
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(10),
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(9),
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(8),
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(7),
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(6),
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(5),
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(4),
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(3),
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(2),
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(1),
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(0),
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q
,
      ALUMODE(0) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_extra_digit_subtract_del_opt_has_pipe_first_q
,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 15),
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 14),
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 13),
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 12),
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 11),
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 10),
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 9),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 8),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 7),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 6),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 5),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 4),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 3),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digit_op(2, 2),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(33),
      P(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(32),
      P(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(31),
      P(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(30),
      P(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(29),
      P(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(28),
      P(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(27),
      P(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(26),
      P(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(25),
      P(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(24),
      P(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(23),
      P(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(22),
      P(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(21),
      P(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(20),
      P(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(19),
      P(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(18),
      P(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(17),
      P(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(16),
      P(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(15),
      P(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(14),
      P(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(13),
      P(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(12),
      P(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(11),
      P(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(10),
      P(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(9),
      P(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(8),
      P(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(7),
      P(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(6),
      P(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(5),
      P(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(4),
      P(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(3),
      P(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(2),
      P(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(1),
      P(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_out_ed(0),
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(18),
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(17),
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(16),
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(15),
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(14),
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(13),
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(12),
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(11),
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(10),
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(9),
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(8),
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(7),
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(6),
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(5),
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(4),
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(3),
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(2),
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_estimate_d(1),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      PCOUT(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_47_UNCONNECTED
,
      PCOUT(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_46_UNCONNECTED
,
      PCOUT(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_45_UNCONNECTED
,
      PCOUT(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_44_UNCONNECTED
,
      PCOUT(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_43_UNCONNECTED
,
      PCOUT(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_42_UNCONNECTED
,
      PCOUT(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_41_UNCONNECTED
,
      PCOUT(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_40_UNCONNECTED
,
      PCOUT(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_39_UNCONNECTED
,
      PCOUT(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_38_UNCONNECTED
,
      PCOUT(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_37_UNCONNECTED
,
      PCOUT(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_36_UNCONNECTED
,
      PCOUT(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_35_UNCONNECTED
,
      PCOUT(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_34_UNCONNECTED
,
      PCOUT(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_33_UNCONNECTED
,
      PCOUT(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_32_UNCONNECTED
,
      PCOUT(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_31_UNCONNECTED
,
      PCOUT(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_30_UNCONNECTED
,
      PCOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_29_UNCONNECTED
,
      PCOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_28_UNCONNECTED
,
      PCOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_27_UNCONNECTED
,
      PCOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_26_UNCONNECTED
,
      PCOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_25_UNCONNECTED
,
      PCOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_24_UNCONNECTED
,
      PCOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_23_UNCONNECTED
,
      PCOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_22_UNCONNECTED
,
      PCOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_21_UNCONNECTED
,
      PCOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_20_UNCONNECTED
,
      PCOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_19_UNCONNECTED
,
      PCOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_18_UNCONNECTED
,
      PCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_17_UNCONNECTED
,
      PCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_16_UNCONNECTED
,
      PCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_15_UNCONNECTED
,
      PCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_14_UNCONNECTED
,
      PCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_13_UNCONNECTED
,
      PCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_12_UNCONNECTED
,
      PCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_11_UNCONNECTED
,
      PCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_10_UNCONNECTED
,
      PCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_9_UNCONNECTED
,
      PCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_8_UNCONNECTED
,
      PCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_7_UNCONNECTED
,
      PCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_6_UNCONNECTED
,
      PCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_5_UNCONNECTED
,
      PCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_4_UNCONNECTED
,
      PCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_3_UNCONNECTED
,
      PCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_2_UNCONNECTED
,
      PCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_1_UNCONNECTED
,
      PCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_multadd_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PCOUT_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(31) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(17),
      C(30) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(16),
      C(29) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(15),
      C(28) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(14),
      C(27) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(13),
      C(26) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(12),
      C(25) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(11),
      C(24) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(10),
      C(23) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(9),
      C(22) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(8),
      C(21) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(7),
      C(20) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(6),
      C(19) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(5),
      C(18) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(4),
      C(17) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(3),
      C(16) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(2),
      C(15) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(1),
      C(14) => 
U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_digits_carrysave_d(0),
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(14),
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(13),
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(12),
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(11),
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(10),
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(9),
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(8),
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(7),
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(6),
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(5),
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(4),
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(3),
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(2),
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_extra_pp_digit_op(1),
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCOUT(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(47),
      PCOUT(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(46),
      PCOUT(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(45),
      PCOUT(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(44),
      PCOUT(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(43),
      PCOUT(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(42),
      PCOUT(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(41),
      PCOUT(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(40),
      PCOUT(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(39),
      PCOUT(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(38),
      PCOUT(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(37),
      PCOUT(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(36),
      PCOUT(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(35),
      PCOUT(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(34),
      PCOUT(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(33),
      PCOUT(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(32),
      PCOUT(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(31),
      PCOUT(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(30),
      PCOUT(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(29),
      PCOUT(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(28),
      PCOUT(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(27),
      PCOUT(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(26),
      PCOUT(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(25),
      PCOUT(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(24),
      PCOUT(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(23),
      PCOUT(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(22),
      PCOUT(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(21),
      PCOUT(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(20),
      PCOUT(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(19),
      PCOUT(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(18),
      PCOUT(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(17),
      PCOUT(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(16),
      PCOUT(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(15),
      PCOUT(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(14),
      PCOUT(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(13),
      PCOUT(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(12),
      PCOUT(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(11),
      PCOUT(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(10),
      PCOUT(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(9),
      PCOUT(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(8),
      PCOUT(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(7),
      PCOUT(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(6),
      PCOUT(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(5),
      PCOUT(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(4),
      PCOUT(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(3),
      PCOUT(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(2),
      PCOUT(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(1),
      PCOUT(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_p_extra_casc(0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED
,
      P(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED
,
      P(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED
,
      P(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED
,
      P(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED
,
      P(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED
,
      P(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED
,
      P(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED
,
      P(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED
,
      P(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED
,
      P(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED
,
      P(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_extra_digits_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED
,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 18),
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 17),
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 16),
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 15),
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 14),
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 13),
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 12),
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 11),
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 10),
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 9),
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 8),
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 7),
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 6),
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 5),
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 4),
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 3),
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 2),
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 1),
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(0, 0),
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCOUT(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 47),
      PCOUT(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 46),
      PCOUT(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 45),
      PCOUT(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 44),
      PCOUT(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 43),
      PCOUT(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 42),
      PCOUT(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 41),
      PCOUT(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 40),
      PCOUT(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 39),
      PCOUT(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 38),
      PCOUT(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 37),
      PCOUT(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 36),
      PCOUT(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 35),
      PCOUT(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 34),
      PCOUT(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 33),
      PCOUT(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 32),
      PCOUT(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 31),
      PCOUT(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 30),
      PCOUT(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 29),
      PCOUT(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 28),
      PCOUT(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 27),
      PCOUT(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 26),
      PCOUT(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 25),
      PCOUT(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 24),
      PCOUT(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 23),
      PCOUT(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 22),
      PCOUT(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 21),
      PCOUT(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 20),
      PCOUT(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 19),
      PCOUT(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 18),
      PCOUT(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 17),
      PCOUT(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 16),
      PCOUT(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 15),
      PCOUT(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 14),
      PCOUT(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 13),
      PCOUT(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 12),
      PCOUT(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 11),
      PCOUT(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 10),
      PCOUT(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 9),
      PCOUT(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 8),
      PCOUT(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 7),
      PCOUT(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 6),
      PCOUT(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 5),
      PCOUT(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 4),
      PCOUT(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 3),
      PCOUT(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 2),
      PCOUT(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 1),
      PCOUT(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(0, 0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED
,
      P(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED
,
      P(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED
,
      P(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED
,
      P(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED
,
      P(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED
,
      P(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED
,
      P(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED
,
      P(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED
,
      P(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED
,
      P(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED
,
      P(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_0_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 18),
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 17),
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 16),
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 15),
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 14),
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 13),
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 12),
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 11),
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 10),
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 9),
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 8),
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 7),
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 6),
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 5),
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 4),
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 3),
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 2),
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 1),
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(1, 0),
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_17_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_15_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_14_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_13_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_12_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_11_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_10_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_9_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_8_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_7_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_6_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_5_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_4_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_3_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_2_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_1_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_32_Q,
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_31_Q,
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_30_Q,
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_29_Q,
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_28_Q,
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_27_Q,
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_26_Q,
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_25_Q,
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_24_Q,
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_23_Q,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_22_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_21_Q,
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_20_Q,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_19_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_1_18_Q,
      PCOUT(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 47),
      PCOUT(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 46),
      PCOUT(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 45),
      PCOUT(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 44),
      PCOUT(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 43),
      PCOUT(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 42),
      PCOUT(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 41),
      PCOUT(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 40),
      PCOUT(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 39),
      PCOUT(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 38),
      PCOUT(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 37),
      PCOUT(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 36),
      PCOUT(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 35),
      PCOUT(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 34),
      PCOUT(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 33),
      PCOUT(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 32),
      PCOUT(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 31),
      PCOUT(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 30),
      PCOUT(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 29),
      PCOUT(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 28),
      PCOUT(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 27),
      PCOUT(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 26),
      PCOUT(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 25),
      PCOUT(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 24),
      PCOUT(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 23),
      PCOUT(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 22),
      PCOUT(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 21),
      PCOUT(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 20),
      PCOUT(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 19),
      PCOUT(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 18),
      PCOUT(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 17),
      PCOUT(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 16),
      PCOUT(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 15),
      PCOUT(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 14),
      PCOUT(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 13),
      PCOUT(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 12),
      PCOUT(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 11),
      PCOUT(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 10),
      PCOUT(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 9),
      PCOUT(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 8),
      PCOUT(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 7),
      PCOUT(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 6),
      PCOUT(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 5),
      PCOUT(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 4),
      PCOUT(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 3),
      PCOUT(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 2),
      PCOUT(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 1),
      PCOUT(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(1, 0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED
,
      P(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED
,
      P(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED
,
      P(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED
,
      P(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED
,
      P(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED
,
      P(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED
,
      P(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED
,
      P(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED
,
      P(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED
,
      P(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED
,
      P(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_1_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive : 
DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 1,
      CREG => 1,
      MASK => X"3FFFFFFFFFFF",
      MREG => 0,
      MULTCARRYINREG => 0,
      OPMODEREG => 1,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "NONE",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CECTRL => aclken,
      CLK => aclk,
      PATTERNBDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNBDETECT_UNCONNECTED
,
      RSTC => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_MULTSIGNOUT_UNCONNECTED
,
      CEC => aclken,
      RSTM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      MULTSIGNIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEB2 => aclken,
      RSTCTRL => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEP => aclken,
      CARRYCASCOUT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYCASCOUT_UNCONNECTED
,
      RSTA => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CECARRYIN => aclken,
      UNDERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_UNDERFLOW_UNCONNECTED
,
      PATTERNDETECT => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_PATTERNDETECT_UNCONNECTED
,
      RSTALUMODE => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTALLCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEALUMODE => aclken,
      CEA2 => aclken,
      CEA1 => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTB => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CEMULTCARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OVERFLOW => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_OVERFLOW_UNCONNECTED
,
      CEM => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYCASCIN => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      RSTP => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYINSEL(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(5) => N0,
      OPMODE(4) => N0,
      OPMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      OPMODE(1) => N0,
      OPMODE(0) => N0,
      C(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 18),
      C(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 17),
      C(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 16),
      C(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 15),
      C(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 14),
      C(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 13),
      C(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 12),
      C(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 11),
      C(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 10),
      C(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 9),
      C(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 8),
      C(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 7),
      C(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 6),
      C(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 5),
      C(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 4),
      C(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 3),
      C(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 2),
      C(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 1),
      C(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_carrysave(2, 0),
      C(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      C(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      B(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_17_Q,
      B(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_16_Q,
      B(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_15_Q,
      B(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_14_Q,
      B(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_13_Q,
      B(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_12_Q,
      B(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_11_Q,
      B(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_10_Q,
      B(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_9_Q,
      B(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_8_Q,
      B(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_7_Q,
      B(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_6_Q,
      B(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_5_Q,
      B(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_4_Q,
      B(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_3_Q,
      B(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_2_Q,
      B(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_1_Q,
      B(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_0_Q,
      A(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_47_Q,
      A(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_46_Q,
      A(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_45_Q,
      A(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_44_Q,
      A(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_43_Q,
      A(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_42_Q,
      A(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_41_Q,
      A(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_40_Q,
      A(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_39_Q,
      A(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_38_Q,
      A(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_37_Q,
      A(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_36_Q,
      A(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_35_Q,
      A(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_34_Q,
      A(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_33_Q,
      A(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_32_Q,
      A(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_31_Q,
      A(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_30_Q,
      A(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_29_Q,
      A(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_28_Q,
      A(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_27_Q,
      A(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_26_Q,
      A(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_25_Q,
      A(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_24_Q,
      A(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_23_Q,
      A(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_22_Q,
      A(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_21_Q,
      A(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_20_Q,
      A(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_19_Q,
      A(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_2_18_Q,
      PCOUT(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 47),
      PCOUT(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 46),
      PCOUT(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 45),
      PCOUT(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 44),
      PCOUT(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 43),
      PCOUT(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 42),
      PCOUT(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 41),
      PCOUT(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 40),
      PCOUT(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 39),
      PCOUT(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 38),
      PCOUT(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 37),
      PCOUT(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 36),
      PCOUT(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 35),
      PCOUT(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 34),
      PCOUT(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 33),
      PCOUT(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 32),
      PCOUT(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 31),
      PCOUT(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 30),
      PCOUT(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 29),
      PCOUT(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 28),
      PCOUT(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 27),
      PCOUT(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 26),
      PCOUT(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 25),
      PCOUT(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 24),
      PCOUT(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 23),
      PCOUT(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 22),
      PCOUT(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 21),
      PCOUT(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 20),
      PCOUT(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 19),
      PCOUT(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 18),
      PCOUT(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 17),
      PCOUT(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 16),
      PCOUT(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 15),
      PCOUT(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 14),
      PCOUT(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 13),
      PCOUT(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 12),
      PCOUT(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 11),
      PCOUT(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 10),
      PCOUT(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 9),
      PCOUT(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 8),
      PCOUT(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 7),
      PCOUT(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 6),
      PCOUT(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 5),
      PCOUT(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 4),
      PCOUT(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 3),
      PCOUT(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 2),
      PCOUT(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 1),
      PCOUT(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_p_casc(2, 0),
      ACOUT(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_29_UNCONNECTED
,
      ACOUT(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_28_UNCONNECTED
,
      ACOUT(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_27_UNCONNECTED
,
      ACOUT(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_26_UNCONNECTED
,
      ACOUT(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_25_UNCONNECTED
,
      ACOUT(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_24_UNCONNECTED
,
      ACOUT(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_23_UNCONNECTED
,
      ACOUT(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_22_UNCONNECTED
,
      ACOUT(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_21_UNCONNECTED
,
      ACOUT(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_20_UNCONNECTED
,
      ACOUT(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_19_UNCONNECTED
,
      ACOUT(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_18_UNCONNECTED
,
      ACOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_17_UNCONNECTED
,
      ACOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_16_UNCONNECTED
,
      ACOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_15_UNCONNECTED
,
      ACOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_14_UNCONNECTED
,
      ACOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_13_UNCONNECTED
,
      ACOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_12_UNCONNECTED
,
      ACOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_11_UNCONNECTED
,
      ACOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_10_UNCONNECTED
,
      ACOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_9_UNCONNECTED
,
      ACOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_8_UNCONNECTED
,
      ACOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_7_UNCONNECTED
,
      ACOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_6_UNCONNECTED
,
      ACOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_5_UNCONNECTED
,
      ACOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_4_UNCONNECTED
,
      ACOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_3_UNCONNECTED
,
      ACOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_2_UNCONNECTED
,
      ACOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_1_UNCONNECTED
,
      ACOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_ACOUT_0_UNCONNECTED
,
      PCIN(47) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(46) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(45) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(44) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(43) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(42) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(41) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(40) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(39) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(38) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(37) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(36) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(35) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(34) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(33) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(32) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(31) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(30) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      PCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ALUMODE(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      CARRYOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_3_UNCONNECTED
,
      CARRYOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_2_UNCONNECTED
,
      CARRYOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_1_UNCONNECTED
,
      CARRYOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_CARRYOUT_0_UNCONNECTED
,
      BCIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      BCOUT(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_17_UNCONNECTED
,
      BCOUT(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_16_UNCONNECTED
,
      BCOUT(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_15_UNCONNECTED
,
      BCOUT(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_14_UNCONNECTED
,
      BCOUT(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_13_UNCONNECTED
,
      BCOUT(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_12_UNCONNECTED
,
      BCOUT(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_11_UNCONNECTED
,
      BCOUT(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_10_UNCONNECTED
,
      BCOUT(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_9_UNCONNECTED
,
      BCOUT(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_8_UNCONNECTED
,
      BCOUT(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_7_UNCONNECTED
,
      BCOUT(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_6_UNCONNECTED
,
      BCOUT(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_5_UNCONNECTED
,
      BCOUT(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_4_UNCONNECTED
,
      BCOUT(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_3_UNCONNECTED
,
      BCOUT(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_2_UNCONNECTED
,
      BCOUT(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_1_UNCONNECTED
,
      BCOUT(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_BCOUT_0_UNCONNECTED
,
      P(47) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_47_UNCONNECTED
,
      P(46) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_46_UNCONNECTED
,
      P(45) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_45_UNCONNECTED
,
      P(44) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_44_UNCONNECTED
,
      P(43) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_43_UNCONNECTED
,
      P(42) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_42_UNCONNECTED
,
      P(41) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_41_UNCONNECTED
,
      P(40) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_40_UNCONNECTED
,
      P(39) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_39_UNCONNECTED
,
      P(38) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_38_UNCONNECTED
,
      P(37) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_37_UNCONNECTED
,
      P(36) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_36_UNCONNECTED
,
      P(35) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_35_UNCONNECTED
,
      P(34) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_34_UNCONNECTED
,
      P(33) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_33_UNCONNECTED
,
      P(32) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_32_UNCONNECTED
,
      P(31) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_31_UNCONNECTED
,
      P(30) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_30_UNCONNECTED
,
      P(29) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_29_UNCONNECTED
,
      P(28) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_28_UNCONNECTED
,
      P(27) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_27_UNCONNECTED
,
      P(26) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_26_UNCONNECTED
,
      P(25) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_25_UNCONNECTED
,
      P(24) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_24_UNCONNECTED
,
      P(23) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_23_UNCONNECTED
,
      P(22) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_22_UNCONNECTED
,
      P(21) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_21_UNCONNECTED
,
      P(20) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_20_UNCONNECTED
,
      P(19) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_19_UNCONNECTED
,
      P(18) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_18_UNCONNECTED
,
      P(17) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_17_UNCONNECTED
,
      P(16) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_16_UNCONNECTED
,
      P(15) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_15_UNCONNECTED
,
      P(14) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_14_UNCONNECTED
,
      P(13) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_13_UNCONNECTED
,
      P(12) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_12_UNCONNECTED
,
      P(11) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_11_UNCONNECTED
,
      P(10) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_10_UNCONNECTED
,
      P(9) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_9_UNCONNECTED
,
      P(8) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_8_UNCONNECTED
,
      P(7) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_7_UNCONNECTED
,
      P(6) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_6_UNCONNECTED
,
      P(5) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_5_UNCONNECTED
,
      P(4) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_4_UNCONNECTED
,
      P(3) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_3_UNCONNECTED
,
      P(2) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_2_UNCONNECTED
,
      P(1) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_1_UNCONNECTED
,
      P(0) => 
NLW_U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_i_splice_2_i_add_i_synth_option_i_synth_model_opt_vx5_i_uniwrap_i_primitive_P_0_UNCONNECTED
,
      ACIN(29) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(28) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(27) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(26) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(25) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(24) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(23) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(22) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(21) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(20) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(19) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(18) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(17) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(16) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(15) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(14) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(13) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(12) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(11) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(10) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(9) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(8) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(7) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(6) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(5) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(4) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(3) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(2) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(1) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q,
      ACIN(0) => U0_i_synth_i_nonzero_fract_i_synth_opt_high_radix_i_nonzero_fract_i_high_radix_i_iterative_unit_abconcat_bus_0_0_Q
    );

end STRUCTURE;

-- synthesis translate_on
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fifo_fg84_26bc5f646d342e7f.vhd when simulating
-- the core, fifo_fg84_26bc5f646d342e7f. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fifo_fg84_26bc5f646d342e7f IS
  PORT (
    clk : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC
  );
END fifo_fg84_26bc5f646d342e7f;

ARCHITECTURE fifo_fg84_26bc5f646d342e7f_a OF fifo_fg84_26bc5f646d342e7f IS
-- synthesis translate_off
COMPONENT wrapped_fifo_fg84_26bc5f646d342e7f
  PORT (
    clk : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(26 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fifo_fg84_26bc5f646d342e7f USE ENTITY XilinxCoreLib.fifo_generator_v8_4(behavioral)
    GENERIC MAP (
      c_add_ngc_constraint => 0,
      c_application_type_axis => 0,
      c_application_type_rach => 0,
      c_application_type_rdch => 0,
      c_application_type_wach => 0,
      c_application_type_wdch => 0,
      c_application_type_wrch => 0,
      c_axi_addr_width => 32,
      c_axi_aruser_width => 1,
      c_axi_awuser_width => 1,
      c_axi_buser_width => 1,
      c_axi_data_width => 64,
      c_axi_id_width => 4,
      c_axi_ruser_width => 1,
      c_axi_type => 0,
      c_axi_wuser_width => 1,
      c_axis_tdata_width => 64,
      c_axis_tdest_width => 4,
      c_axis_tid_width => 8,
      c_axis_tkeep_width => 4,
      c_axis_tstrb_width => 4,
      c_axis_tuser_width => 4,
      c_axis_type => 0,
      c_common_clock => 1,
      c_count_type => 0,
      c_data_count_width => 8,
      c_default_value => "BlankString",
      c_din_width => 27,
      c_din_width_axis => 1,
      c_din_width_rach => 32,
      c_din_width_rdch => 64,
      c_din_width_wach => 32,
      c_din_width_wdch => 64,
      c_din_width_wrch => 2,
      c_dout_rst_val => "0",
      c_dout_width => 27,
      c_enable_rlocs => 0,
      c_enable_rst_sync => 1,
      c_error_injection_type => 0,
      c_error_injection_type_axis => 0,
      c_error_injection_type_rach => 0,
      c_error_injection_type_rdch => 0,
      c_error_injection_type_wach => 0,
      c_error_injection_type_wdch => 0,
      c_error_injection_type_wrch => 0,
      c_family => "virtex6",
      c_full_flags_rst_val => 0,
      c_has_almost_empty => 0,
      c_has_almost_full => 0,
      c_has_axi_aruser => 0,
      c_has_axi_awuser => 0,
      c_has_axi_buser => 0,
      c_has_axi_rd_channel => 0,
      c_has_axi_ruser => 0,
      c_has_axi_wr_channel => 0,
      c_has_axi_wuser => 0,
      c_has_axis_tdata => 0,
      c_has_axis_tdest => 0,
      c_has_axis_tid => 0,
      c_has_axis_tkeep => 0,
      c_has_axis_tlast => 0,
      c_has_axis_tready => 1,
      c_has_axis_tstrb => 0,
      c_has_axis_tuser => 0,
      c_has_backup => 0,
      c_has_data_count => 0,
      c_has_data_counts_axis => 0,
      c_has_data_counts_rach => 0,
      c_has_data_counts_rdch => 0,
      c_has_data_counts_wach => 0,
      c_has_data_counts_wdch => 0,
      c_has_data_counts_wrch => 0,
      c_has_int_clk => 0,
      c_has_master_ce => 0,
      c_has_meminit_file => 0,
      c_has_overflow => 0,
      c_has_prog_flags_axis => 0,
      c_has_prog_flags_rach => 0,
      c_has_prog_flags_rdch => 0,
      c_has_prog_flags_wach => 0,
      c_has_prog_flags_wdch => 0,
      c_has_prog_flags_wrch => 0,
      c_has_rd_data_count => 0,
      c_has_rd_rst => 0,
      c_has_rst => 0,
      c_has_slave_ce => 0,
      c_has_srst => 0,
      c_has_underflow => 0,
      c_has_valid => 0,
      c_has_wr_ack => 0,
      c_has_wr_data_count => 0,
      c_has_wr_rst => 0,
      c_implementation_type => 0,
      c_implementation_type_axis => 1,
      c_implementation_type_rach => 1,
      c_implementation_type_rdch => 1,
      c_implementation_type_wach => 1,
      c_implementation_type_wdch => 1,
      c_implementation_type_wrch => 1,
      c_init_wr_pntr_val => 0,
      c_interface_type => 0,
      c_memory_type => 2,
      c_mif_file_name => "BlankString",
      c_msgon_val => 1,
      c_optimization_mode => 0,
      c_overflow_low => 0,
      c_preload_latency => 0,
      c_preload_regs => 1,
      c_prim_fifo_type => "512x36",
      c_prog_empty_thresh_assert_val => 4,
      c_prog_empty_thresh_assert_val_axis => 1022,
      c_prog_empty_thresh_assert_val_rach => 1022,
      c_prog_empty_thresh_assert_val_rdch => 1022,
      c_prog_empty_thresh_assert_val_wach => 1022,
      c_prog_empty_thresh_assert_val_wdch => 1022,
      c_prog_empty_thresh_assert_val_wrch => 1022,
      c_prog_empty_thresh_negate_val => 5,
      c_prog_empty_type => 0,
      c_prog_empty_type_axis => 5,
      c_prog_empty_type_rach => 5,
      c_prog_empty_type_rdch => 5,
      c_prog_empty_type_wach => 5,
      c_prog_empty_type_wdch => 5,
      c_prog_empty_type_wrch => 5,
      c_prog_full_thresh_assert_val => 127,
      c_prog_full_thresh_assert_val_axis => 1023,
      c_prog_full_thresh_assert_val_rach => 1023,
      c_prog_full_thresh_assert_val_rdch => 1023,
      c_prog_full_thresh_assert_val_wach => 1023,
      c_prog_full_thresh_assert_val_wdch => 1023,
      c_prog_full_thresh_assert_val_wrch => 1023,
      c_prog_full_thresh_negate_val => 126,
      c_prog_full_type => 0,
      c_prog_full_type_axis => 5,
      c_prog_full_type_rach => 5,
      c_prog_full_type_rdch => 5,
      c_prog_full_type_wach => 5,
      c_prog_full_type_wdch => 5,
      c_prog_full_type_wrch => 5,
      c_rach_type => 0,
      c_rd_data_count_width => 8,
      c_rd_depth => 128,
      c_rd_freq => 1,
      c_rd_pntr_width => 7,
      c_rdch_type => 0,
      c_reg_slice_mode_axis => 0,
      c_reg_slice_mode_rach => 0,
      c_reg_slice_mode_rdch => 0,
      c_reg_slice_mode_wach => 0,
      c_reg_slice_mode_wdch => 0,
      c_reg_slice_mode_wrch => 0,
      c_synchronizer_stage => 2,
      c_underflow_low => 0,
      c_use_common_overflow => 0,
      c_use_common_underflow => 0,
      c_use_default_settings => 0,
      c_use_dout_rst => 0,
      c_use_ecc => 0,
      c_use_ecc_axis => 0,
      c_use_ecc_rach => 0,
      c_use_ecc_rdch => 0,
      c_use_ecc_wach => 0,
      c_use_ecc_wdch => 0,
      c_use_ecc_wrch => 0,
      c_use_embedded_reg => 0,
      c_use_fifo16_flags => 0,
      c_use_fwft_data_count => 1,
      c_valid_low => 0,
      c_wach_type => 0,
      c_wdch_type => 0,
      c_wr_ack_low => 0,
      c_wr_data_count_width => 8,
      c_wr_depth => 128,
      c_wr_depth_axis => 1024,
      c_wr_depth_rach => 16,
      c_wr_depth_rdch => 1024,
      c_wr_depth_wach => 16,
      c_wr_depth_wdch => 1024,
      c_wr_depth_wrch => 16,
      c_wr_freq => 1,
      c_wr_pntr_width => 7,
      c_wr_pntr_width_axis => 10,
      c_wr_pntr_width_rach => 4,
      c_wr_pntr_width_rdch => 10,
      c_wr_pntr_width_wach => 4,
      c_wr_pntr_width_wdch => 10,
      c_wr_pntr_width_wrch => 4,
      c_wr_response_latency => 1,
      c_wrch_type => 0
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fifo_fg84_26bc5f646d342e7f
  PORT MAP (
    clk => clk,
    din => din,
    wr_en => wr_en,
    rd_en => rd_en,
    dout => dout,
    full => full,
    empty => empty
  );
-- synthesis translate_on

END fifo_fg84_26bc5f646d342e7f_a;
--------------------------------------------------------------------------------
--     (c) Copyright 1995 - 2010 Xilinx, Inc. All rights reserved.            --
--                                                                            --
--     This file contains confidential and proprietary information            --
--     of Xilinx, Inc. and is protected under U.S. and                        --
--     international copyright and other intellectual property                --
--     laws.                                                                  --
--                                                                            --
--     DISCLAIMER                                                             --
--     This disclaimer is not a license and does not grant any                --
--     rights to the materials distributed herewith. Except as                --
--     otherwise provided in a valid license issued to you by                 --
--     Xilinx, and to the maximum extent permitted by applicable              --
--     law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND                --
--     WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES            --
--     AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING              --
--     BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-                 --
--     INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and               --
--     (2) Xilinx shall not be liable (whether in contract or tort,           --
--     including negligence, or under any other theory of                     --
--     liability) for any loss or damage of any kind or nature                --
--     related to, arising under or in connection with these                  --
--     materials, including for any direct, or any indirect,                  --
--     special, incidental, or consequential loss or damage                   --
--     (including loss of data, profits, goodwill, or any type of             --
--     loss or damage suffered as a result of any action brought              --
--     by a third party) even if such damage or loss was                      --
--     reasonably foreseeable or Xilinx had been advised of the               --
--     possibility of the same.                                               --
--                                                                            --
--     CRITICAL APPLICATIONS                                                  --
--     Xilinx products are not designed or intended to be fail-               --
--     safe, or for use in any application requiring fail-safe                --
--     performance, such as life-support or safety devices or                 --
--     systems, Class III medical devices, nuclear facilities,                --
--     applications related to the deployment of airbags, or any              --
--     other applications that could lead to death, personal                  --
--     injury, or severe property or environmental damage                     --
--     (individually and collectively, "Critical                              --
--     Applications"). Customer assumes the sole risk and                     --
--     liability of any use of Xilinx products in Critical                    --
--     Applications, subject only to applicable laws and                      --
--     regulations governing limitations on product liability.                --
--                                                                            --
--     THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS               --
--     PART OF THIS FILE AT ALL TIMES.                                        --
--------------------------------------------------------------------------------

--  Generated from component ID: xilinx.com:ip:fir_compiler:6.2


-- You must compile the wrapper file fr_cmplr_v6_2_2e31efd348cc2721.vhd when simulating
-- the core, fr_cmplr_v6_2_2e31efd348cc2721. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
Library XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_2_2e31efd348cc2721 IS
	port (
	aclk: in std_logic;
	aclken: in std_logic;
	s_axis_data_tvalid: in std_logic;
	s_axis_data_tready: out std_logic;
	s_axis_data_tdata: in std_logic_vector(47 downto 0);
	m_axis_data_tvalid: out std_logic;
	m_axis_data_tdata: out std_logic_vector(95 downto 0));
END fr_cmplr_v6_2_2e31efd348cc2721;

ARCHITECTURE fr_cmplr_v6_2_2e31efd348cc2721_a OF fr_cmplr_v6_2_2e31efd348cc2721 IS
-- synthesis translate_off
component wrapped_fr_cmplr_v6_2_2e31efd348cc2721
	port (
	aclk: in std_logic;
	aclken: in std_logic;
	s_axis_data_tvalid: in std_logic;
	s_axis_data_tready: out std_logic;
	s_axis_data_tdata: in std_logic_vector(47 downto 0);
	m_axis_data_tvalid: out std_logic;
	m_axis_data_tdata: out std_logic_vector(95 downto 0));
end component;

-- Configuration specification 
	for all : wrapped_fr_cmplr_v6_2_2e31efd348cc2721 use entity XilinxCoreLib.fir_compiler_v6_2(behavioral)
		generic map(
			c_round_mode => 0,
			c_coef_memtype => 2,
			c_has_config_channel => 0,
			c_m_data_has_tready => 0,
			c_col_pipe_len => 4,
			c_coef_reload => 0,
			c_input_rate => 1,
			c_col_config => "14",
			c_coef_mem_packing => 0,
			c_filter_type => 1,
			c_accum_op_path_widths => "45,45",
			c_component_name => "fr_cmplr_v6_2_2e31efd348cc2721",
			c_coef_file => "fr_cmplr_v6_2_2e31efd348cc2721.mif",
			c_reload_tdata_width => 1,
			c_mem_arrangement => 1,
			c_filts_packed => 0,
			c_opbuff_memtype => 0,
			c_num_channels => 1,
			c_data_width => 24,
			c_symmetry => 1,
			c_data_path_src => "0,1",
			c_data_path_sign => "0,0",
			c_config_sync_mode => 0,
			c_latency => 20,
			c_output_rate => 35,
			c_xdevicefamily => "virtex6",
			c_interp_rate => 1,
			c_datapath_memtype => 2,
			c_s_data_tdata_width => 48,
			c_coef_file_lines => 455,
			c_s_data_has_tuser => 0,
			c_s_data_tuser_width => 1,
			c_data_memtype => 0,
			c_output_path_widths => "45,45",
			c_data_path_widths => "24,24",
			c_coef_path_sign => "0,0",
			c_has_aresetn => 0,
			c_decim_rate => 35,
			c_data_has_tlast => 0,
			c_s_data_has_fifo => 0,
			c_oversampling_rate => 1,
			c_channel_pattern => "fixed",
			c_config_packet_size => 0,
			c_coef_path_widths => "16,16",
			c_optimization => 0,
			c_m_data_has_tuser => 0,
			c_num_reload_slots => 1,
			c_coef_path_src => "0,0",
			c_m_data_tdata_width => 96,
			c_has_aclken => 1,
			c_zero_packing_factor => 1,
			c_config_tdata_width => 1,
			c_m_data_tuser_width => 1,
			c_accum_path_widths => "45,45",
			c_num_taps => 841,
			c_ipbuff_memtype => 0,
			c_num_madds => 13,
			c_coef_width => 16,
			c_opt_madds => "none",
			c_num_filts => 1,
			c_data_mem_packing => 0,
			c_ext_mult_cnfg => "none",
			c_output_width => 45,
			c_col_mode => 0);
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_2_2e31efd348cc2721
		port map (
			aclk => aclk,
			aclken => aclken,
			s_axis_data_tvalid => s_axis_data_tvalid,
			s_axis_data_tready => s_axis_data_tready,
			s_axis_data_tdata => s_axis_data_tdata,
			m_axis_data_tvalid => m_axis_data_tvalid,
			m_axis_data_tdata => m_axis_data_tdata);
-- synthesis translate_on

END fr_cmplr_v6_2_2e31efd348cc2721_a;

--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_121326a881aa557e.vhd when simulating
-- the core, fr_cmplr_v6_3_121326a881aa557e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_121326a881aa557e IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END fr_cmplr_v6_3_121326a881aa557e;

ARCHITECTURE fr_cmplr_v6_3_121326a881aa557e_a OF fr_cmplr_v6_3_121326a881aa557e IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_121326a881aa557e
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_121326a881aa557e USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "43",
      c_accum_path_widths => "31,30",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_121326a881aa557e.mif",
      c_coef_file_lines => 42,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0,0",
      c_coef_path_src => "0,0",
      c_coef_path_widths => "16,16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "21",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_121326a881aa557e",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 0,
      c_data_path_sign => "1,0",
      c_data_path_src => "0,1",
      c_data_path_widths => "13,13",
      c_data_width => 26,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "0,1,0,13",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 30,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 48,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 1,
      c_num_filts => 1,
      c_num_madds => 21,
      c_num_reload_slots => 1,
      c_num_taps => 81,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "43",
      c_output_rate => 2,
      c_output_width => 43,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 0,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 0,
      c_s_data_tdata_width => 32,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "virtex6",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_121326a881aa557e
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END fr_cmplr_v6_3_121326a881aa557e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_555df73bebb69ee8.vhd when simulating
-- the core, fr_cmplr_v6_3_555df73bebb69ee8. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_555df73bebb69ee8 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END fr_cmplr_v6_3_555df73bebb69ee8;

ARCHITECTURE fr_cmplr_v6_3_555df73bebb69ee8_a OF fr_cmplr_v6_3_555df73bebb69ee8 IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_555df73bebb69ee8
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_555df73bebb69ee8 USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "42",
      c_accum_path_widths => "30,30",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_555df73bebb69ee8.mif",
      c_coef_file_lines => 42,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0,0",
      c_coef_path_src => "0,0",
      c_coef_path_widths => "16,16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "21",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_555df73bebb69ee8",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 0,
      c_data_path_sign => "1,0",
      c_data_path_src => "0,1",
      c_data_path_widths => "12,13",
      c_data_width => 25,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "0,1,0,12",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 30,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 48,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 1,
      c_num_filts => 1,
      c_num_madds => 21,
      c_num_reload_slots => 1,
      c_num_taps => 81,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "42",
      c_output_rate => 2,
      c_output_width => 42,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 0,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 0,
      c_s_data_tdata_width => 32,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "virtex6",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_555df73bebb69ee8
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END fr_cmplr_v6_3_555df73bebb69ee8_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_85eb797d79431254.vhd when simulating
-- the core, fr_cmplr_v6_3_85eb797d79431254. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_85eb797d79431254 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END fr_cmplr_v6_3_85eb797d79431254;

ARCHITECTURE fr_cmplr_v6_3_85eb797d79431254_a OF fr_cmplr_v6_3_85eb797d79431254 IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_85eb797d79431254
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_85eb797d79431254 USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "41",
      c_accum_path_widths => "41",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_85eb797d79431254.mif",
      c_coef_file_lines => 10,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "5",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_85eb797d79431254",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 0,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "24",
      c_data_width => 24,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 12,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 48,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 1,
      c_num_filts => 1,
      c_num_madds => 5,
      c_num_reload_slots => 1,
      c_num_taps => 17,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "41",
      c_output_rate => 2,
      c_output_width => 41,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 0,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 0,
      c_s_data_tdata_width => 24,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "virtex6",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_85eb797d79431254
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END fr_cmplr_v6_3_85eb797d79431254_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_8dca82a218dd87c6.vhd when simulating
-- the core, fr_cmplr_v6_3_8dca82a218dd87c6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_8dca82a218dd87c6 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(39 DOWNTO 0)
  );
END fr_cmplr_v6_3_8dca82a218dd87c6;

ARCHITECTURE fr_cmplr_v6_3_8dca82a218dd87c6_a OF fr_cmplr_v6_3_8dca82a218dd87c6 IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_8dca82a218dd87c6
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(39 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_8dca82a218dd87c6 USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "34",
      c_accum_path_widths => "34",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_8dca82a218dd87c6.mif",
      c_coef_file_lines => 29,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "29",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_8dca82a218dd87c6",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 0,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "16",
      c_data_width => 16,
      c_datapath_memtype => 0,
      c_decim_rate => 1,
      c_ext_mult_cnfg => "none",
      c_filter_type => 0,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 35,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 40,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 1,
      c_num_filts => 1,
      c_num_madds => 29,
      c_num_reload_slots => 1,
      c_num_taps => 57,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "34",
      c_output_rate => 1,
      c_output_width => 34,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 0,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 0,
      c_s_data_tdata_width => 16,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "virtex6",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_8dca82a218dd87c6
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END fr_cmplr_v6_3_8dca82a218dd87c6_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_8f63af671437d2cb.vhd when simulating
-- the core, fr_cmplr_v6_3_8f63af671437d2cb. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_8f63af671437d2cb IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END fr_cmplr_v6_3_8f63af671437d2cb;

ARCHITECTURE fr_cmplr_v6_3_8f63af671437d2cb_a OF fr_cmplr_v6_3_8f63af671437d2cb IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_8f63af671437d2cb
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_8f63af671437d2cb USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "41",
      c_accum_path_widths => "41",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_8f63af671437d2cb.mif",
      c_coef_file_lines => 10,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "5",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_8f63af671437d2cb",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 0,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "24",
      c_data_width => 24,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 12,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 0,
      c_m_data_tdata_width => 48,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 1,
      c_num_filts => 1,
      c_num_madds => 5,
      c_num_reload_slots => 1,
      c_num_taps => 17,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "41",
      c_output_rate => 2,
      c_output_width => 41,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 0,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 0,
      c_s_data_tdata_width => 24,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "virtex6",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_8f63af671437d2cb
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tdata => m_axis_data_tdata
  );
-- synthesis translate_on

END fr_cmplr_v6_3_8f63af671437d2cb_a;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlclockenablegenerator is
  generic (
    period: integer := 2;
    log_2_period: integer := 0;
    pipeline_regs: integer := 5
  );
  port (
    clk: in std_logic;
    clr: in std_logic;
    ce: out std_logic
  );
end xlclockenablegenerator;
architecture behavior of xlclockenablegenerator is
  component synth_reg_w_init
    generic (
      width: integer;
      init_index: integer;
      init_value: bit_vector;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function size_of_uint(inp: integer; power_of_2: boolean)
    return integer
  is
    constant inp_vec: std_logic_vector(31 downto 0) :=
      integer_to_std_logic_vector(inp,32, xlUnsigned);
    variable result: integer;
  begin
    result := 32;
    for i in 0 to 31 loop
      if inp_vec(i) = '1' then
        result := i;
      end if;
    end loop;
    if power_of_2 then
      return result;
    else
      return result+1;
    end if;
  end;
  function is_power_of_2(inp: std_logic_vector)
    return boolean
  is
    constant width: integer := inp'length;
    variable vec: std_logic_vector(width - 1 downto 0);
    variable single_bit_set: boolean;
    variable more_than_one_bit_set: boolean;
    variable result: boolean;
  begin
    vec := inp;
    single_bit_set := false;
    more_than_one_bit_set := false;
    -- synopsys translate_off
    if (is_XorU(vec)) then
      return false;
    end if;
     -- synopsys translate_on
    if width > 0 then
      for i in 0 to width - 1 loop
        if vec(i) = '1' then
          if single_bit_set then
            more_than_one_bit_set := true;
          end if;
          single_bit_set := true;
        end if;
      end loop;
    end if;
    if (single_bit_set and not(more_than_one_bit_set)) then
      result := true;
    else
      result := false;
    end if;
    return result;
  end;
  function ce_reg_init_val(index, period : integer)
    return integer
  is
     variable result: integer;
   begin
      result := 0;
      if ((index mod period) = 0) then
          result := 1;
      end if;
      return result;
  end;
  function remaining_pipe_regs(num_pipeline_regs, period : integer)
    return integer
  is
     variable factor, result: integer;
  begin
      factor := (num_pipeline_regs / period);
      result := num_pipeline_regs - (period * factor) + 1;
      return result;
  end;

  function sg_min(L, R: INTEGER) return INTEGER is
  begin
      if L < R then
            return L;
      else
            return R;
      end if;
  end;
  constant max_pipeline_regs : integer := 8;
  constant pipe_regs : integer := 5;
  constant num_pipeline_regs : integer := sg_min(pipeline_regs, max_pipeline_regs);
  constant rem_pipeline_regs : integer := remaining_pipe_regs(num_pipeline_regs,period);
  constant period_floor: integer := max(2, period);
  constant power_of_2_counter: boolean :=
    is_power_of_2(integer_to_std_logic_vector(period_floor,32, xlUnsigned));
  constant cnt_width: integer :=
    size_of_uint(period_floor, power_of_2_counter);
  constant clk_for_ce_pulse_minus1: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector((period_floor - 2),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus2: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - 3),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus_regs: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - rem_pipeline_regs),cnt_width, xlUnsigned);
  signal clk_num: unsigned(cnt_width - 1 downto 0) := (others => '0');
  signal ce_vec : std_logic_vector(num_pipeline_regs downto 0);
  signal internal_ce: std_logic_vector(0 downto 0);
  signal cnt_clr, cnt_clr_dly: std_logic_vector (0 downto 0);
begin
  cntr_gen: process(clk)
  begin
    if clk'event and clk = '1'  then
        if ((cnt_clr_dly(0) = '1') or (clr = '1')) then
          clk_num <= (others => '0');
        else
          clk_num <= clk_num + 1;
        end if;
    end if;
  end process;
  clr_gen: process(clk_num, clr)
  begin
    if power_of_2_counter then
      cnt_clr(0) <= clr;
    else
      if (unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus1
          or clr = '1') then
        cnt_clr(0) <= '1';
      else
        cnt_clr(0) <= '0';
      end if;
    end if;
  end process;
  clr_reg: synth_reg_w_init
    generic map (
      width => 1,
      init_index => 0,
      init_value => b"0000",
      latency => 1
    )
    port map (
      i => cnt_clr,
      ce => '1',
      clr => clr,
      clk => clk,
      o => cnt_clr_dly
    );
  pipelined_ce : if period > 1 generate
      ce_gen: process(clk_num)
      begin
          if unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus_regs then
              ce_vec(num_pipeline_regs) <= '1';
          else
              ce_vec(num_pipeline_regs) <= '0';
          end if;
      end process;
      ce_pipeline: for index in num_pipeline_regs downto 1 generate
          ce_reg : synth_reg_w_init
              generic map (
                  width => 1,
                  init_index => ce_reg_init_val(index, period),
                  init_value => b"0000",
                  latency => 1
                  )
              port map (
                  i => ce_vec(index downto index),
                  ce => '1',
                  clr => clr,
                  clk => clk,
                  o => ce_vec(index-1 downto index-1)
                  );
      end generate;
      internal_ce <= ce_vec(0 downto 0);
  end generate;
  generate_clock_enable: if period > 1 generate
    ce <= internal_ce(0);
  end generate;
  generate_clock_enable_constant: if period = 1 generate
    ce <= '1';
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_31a4235b32 is
  port (
    input_port : in std_logic_vector((25 - 1) downto 0);
    output_port : out std_logic_vector((25 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_31a4235b32;


architecture behavior of reinterpret_31a4235b32 is
  signal input_port_1_40: signed((25 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcic_compiler_bb7d6f586f04abec4d028ced88abc8ae is 
  port(
    ce:in std_logic;
    ce_1113:in std_logic;
    ce_logic_1:in std_logic;
    clk:in std_logic;
    clk_1113:in std_logic;
    clk_logic_1:in std_logic;
    m_axis_data_tdata_data:out std_logic_vector(24 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_data:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic
  );
end xlcic_compiler_bb7d6f586f04abec4d028ced88abc8ae;


architecture behavior of xlcic_compiler_bb7d6f586f04abec4d028ced88abc8ae  is
  component cc_cmplr_v3_0_75f3b28f5ac4aa5e
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_captured: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_or_captured_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_data_ps_net <= m_axis_data_tdata_net(24 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_data;
  m_axis_data_tdata_data_ps_net_or_captured_net <= m_axis_data_tdata_data_ps_net or m_axis_data_tdata_data_ps_net_captured;
m_axis_data_tdata_data_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net_or_captured_net,
        ce => ce_1113,
        clr => '0',
        clk => clk_1113, 
        o => m_axis_data_tdata_data
    );
m_axis_data_tdata_data_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1113, 
        o => m_axis_data_tdata_data_ps_net_captured
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_1113,
        clr => '0',
        clk => clk_1113, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1113, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  cc_cmplr_v3_0_75f3b28f5ac4aa5e_instance : cc_cmplr_v3_0_75f3b28f5ac4aa5e
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_1
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcordic_c062cc3a2d77ede2032de397150e15cd is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_phase:out std_logic_vector(24 downto 0);
    m_axis_dout_tdata_real:out std_logic_vector(24 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_cartesian_tdata_imag:in std_logic_vector(24 downto 0);
    s_axis_cartesian_tdata_real:in std_logic_vector(24 downto 0);
    s_axis_cartesian_tvalid:in std_logic
  );
end xlcordic_c062cc3a2d77ede2032de397150e15cd;


architecture behavior of xlcordic_c062cc3a2d77ede2032de397150e15cd  is
  component crdc_v5_0_ac582be577bf89c0
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(63 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_cartesian_tdata:in std_logic_vector(63 downto 0);
      s_axis_cartesian_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
signal s_axis_cartesian_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_phase <= m_axis_dout_tdata_net(56 downto 32);
  m_axis_dout_tdata_real <= m_axis_dout_tdata_net(24 downto 0);
  s_axis_cartesian_tdata_net(56 downto 32) <= s_axis_cartesian_tdata_imag;
  s_axis_cartesian_tdata_net(24 downto 0) <= s_axis_cartesian_tdata_real;
  crdc_v5_0_ac582be577bf89c0_instance : crdc_v5_0_ac582be577bf89c0
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_cartesian_tdata=>s_axis_cartesian_tdata_net,
      s_axis_cartesian_tvalid=>s_axis_cartesian_tvalid
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcomplex_multiplier_a3a52a268f0fdc1111e428e7f4c7c82c is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_imag:out std_logic_vector(23 downto 0);
    m_axis_dout_tdata_real:out std_logic_vector(23 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_a_tdata_imag:in std_logic_vector(23 downto 0);
    s_axis_a_tdata_real:in std_logic_vector(23 downto 0);
    s_axis_a_tvalid:in std_logic;
    s_axis_b_tdata_imag:in std_logic_vector(23 downto 0);
    s_axis_b_tdata_real:in std_logic_vector(23 downto 0);
    s_axis_b_tvalid:in std_logic
  );
end xlcomplex_multiplier_a3a52a268f0fdc1111e428e7f4c7c82c;


architecture behavior of xlcomplex_multiplier_a3a52a268f0fdc1111e428e7f4c7c82c  is
  component cmpy_v5_0_3b811ae68acefe54
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(47 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_a_tdata:in std_logic_vector(47 downto 0);
      s_axis_a_tvalid:in std_logic;
      s_axis_b_tdata:in std_logic_vector(47 downto 0);
      s_axis_b_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal s_axis_a_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal s_axis_b_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_imag <= m_axis_dout_tdata_net(47 downto 24);
  m_axis_dout_tdata_real <= m_axis_dout_tdata_net(23 downto 0);
  s_axis_a_tdata_net(47 downto 24) <= s_axis_a_tdata_imag;
  s_axis_a_tdata_net(23 downto 0) <= s_axis_a_tdata_real;
  s_axis_b_tdata_net(47 downto 24) <= s_axis_b_tdata_imag;
  s_axis_b_tdata_net(23 downto 0) <= s_axis_b_tdata_real;
  cmpy_v5_0_3b811ae68acefe54_instance : cmpy_v5_0_3b811ae68acefe54
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_a_tdata=>s_axis_a_tdata_net,
      s_axis_a_tvalid=>s_axis_a_tvalid,
      s_axis_b_tdata=>s_axis_b_tdata_net,
      s_axis_b_tvalid=>s_axis_b_tvalid
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_961b43f67a is
  port (
    d : in std_logic_vector((24 - 1) downto 0);
    q : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_961b43f67a;


architecture behavior of delay_961b43f67a is
  signal d_1_22: std_logic_vector((24 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer :=  0;
           reset        : integer :=  0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        rst     : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if ((reg_retiming = 0) and (reset = 0)) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if ((reg_retiming = 1) or (reset = 1)) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => rst,
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_b62f4240f0 is
  port (
    input_port : in std_logic_vector((24 - 1) downto 0);
    output_port : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_b62f4240f0;


architecture behavior of reinterpret_b62f4240f0 is
  signal input_port_1_40: signed((24 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_db690cb1dac026c47ff98d5afcede74f is 
  port(
    ce:in std_logic;
    ce_logic_1:in std_logic;
    clk:in std_logic;
    clk_logic_1:in std_logic;
    m_axis_data_tdata:out std_logic_vector(33 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(15 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_db690cb1dac026c47ff98d5afcede74f;


architecture behavior of xlfir_compiler_db690cb1dac026c47ff98d5afcede74f  is
  component fr_cmplr_v6_3_8dca82a218dd87c6
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(39 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(15 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(39 downto 0) := (others=>'0');
signal s_axis_data_tdata_net: std_logic_vector(15 downto 0) := (others=>'0');
begin
  m_axis_data_tdata <= m_axis_data_tdata_net(33 downto 0);
  s_axis_data_tdata_net(15 downto 0) <= s_axis_data_tdata;
  fr_cmplr_v6_3_8dca82a218dd87c6_instance : fr_cmplr_v6_3_8dca82a218dd87c6
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_1
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_f394f3309c is
  port (
    op : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_f394f3309c;


architecture behavior of constant_f394f3309c is
begin
  op <= "000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_6d27a36d02c91c0ddc9d14d956c5aca1 is 
  port(
    ce:in std_logic;
    ce_35:in std_logic;
    ce_logic_1:in std_logic;
    clk:in std_logic;
    clk_35:in std_logic;
    clk_logic_1:in std_logic;
    m_axis_data_tdata_path0:out std_logic_vector(44 downto 0);
    m_axis_data_tdata_path1:out std_logic_vector(44 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_path0:in std_logic_vector(23 downto 0);
    s_axis_data_tdata_path1:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_6d27a36d02c91c0ddc9d14d956c5aca1;


architecture behavior of xlfir_compiler_6d27a36d02c91c0ddc9d14d956c5aca1  is
  component fr_cmplr_v6_2_2e31efd348cc2721
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(95 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(47 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(95 downto 0) := (others=>'0');
signal m_axis_data_tdata_path1_ps_net: std_logic_vector(44 downto 0) := (others=>'0');
signal m_axis_data_tdata_path0_ps_net: std_logic_vector(44 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_path1_ps_net <= m_axis_data_tdata_net(92 downto 48);
  m_axis_data_tdata_path0_ps_net <= m_axis_data_tdata_net(44 downto 0);
  s_axis_data_tdata_net(47 downto 24) <= s_axis_data_tdata_path1;
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_path0;
  m_axis_data_tdata_path1_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 45,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_path1_ps_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35, 
        o => m_axis_data_tdata_path1
    );
  m_axis_data_tdata_path0_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 45,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_path0_ps_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35, 
        o => m_axis_data_tdata_path0
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_35, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_2_2e31efd348cc2721_instance : fr_cmplr_v6_2_2e31efd348cc2721
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_1
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_82c3c799ff is
  port (
    input_port : in std_logic_vector((45 - 1) downto 0);
    output_port : out std_logic_vector((45 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_82c3c799ff;


architecture behavior of reinterpret_82c3c799ff is
  signal input_port_1_40: signed((45 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_63d9ad3400f500cbd021770c26f451ad is 
  port(
    ce:in std_logic;
    ce_2782500:in std_logic;
    ce_5565000:in std_logic;
    ce_logic_2782500:in std_logic;
    clk:in std_logic;
    clk_2782500:in std_logic;
    clk_5565000:in std_logic;
    clk_logic_2782500:in std_logic;
    m_axis_data_tdata:out std_logic_vector(40 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_63d9ad3400f500cbd021770c26f451ad;


architecture behavior of xlfir_compiler_63d9ad3400f500cbd021770c26f451ad  is
  component fr_cmplr_v6_3_8f63af671437d2cb
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(47 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(40 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(40 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 41,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_5565000,
        clr => '0',
        clk => clk_5565000, 
        o => m_axis_data_tdata
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_5565000,
        clr => '0',
        clk => clk_5565000, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_5565000, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_8f63af671437d2cb_instance : fr_cmplr_v6_3_8f63af671437d2cb
    port map(
      aclk=>clk,
      aclken=>ce_2782500,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_2782500
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcic_compiler_95547d442151284e81277c01e1dd33ef is 
  port(
    ce:in std_logic;
    ce_1113:in std_logic;
    ce_2782500:in std_logic;
    ce_logic_1113:in std_logic;
    clk:in std_logic;
    clk_1113:in std_logic;
    clk_2782500:in std_logic;
    clk_logic_1113:in std_logic;
    m_axis_data_tdata_data:out std_logic_vector(23 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_data:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic
  );
end xlcic_compiler_95547d442151284e81277c01e1dd33ef;


architecture behavior of xlcic_compiler_95547d442151284e81277c01e1dd33ef  is
  component cc_cmplr_v3_0_2d327f6921329141
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(23 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net: std_logic_vector(23 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_captured: std_logic_vector(23 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_or_captured_net: std_logic_vector(23 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_data_ps_net <= m_axis_data_tdata_net(23 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_data;
  m_axis_data_tdata_data_ps_net_or_captured_net <= m_axis_data_tdata_data_ps_net or m_axis_data_tdata_data_ps_net_captured;
m_axis_data_tdata_data_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 24,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net_or_captured_net,
        ce => ce_2782500,
        clr => '0',
        clk => clk_2782500, 
        o => m_axis_data_tdata_data
    );
m_axis_data_tdata_data_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 24,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_2782500, 
        o => m_axis_data_tdata_data_ps_net_captured
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_2782500,
        clr => '0',
        clk => clk_2782500, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_2782500, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  cc_cmplr_v3_0_2d327f6921329141_instance : cc_cmplr_v3_0_2d327f6921329141
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_1113
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_d0050991ffa08d9151315827675f900b is 
  port(
    ce:in std_logic;
    ce_11130000:in std_logic;
    ce_5565000:in std_logic;
    ce_logic_5565000:in std_logic;
    clk:in std_logic;
    clk_11130000:in std_logic;
    clk_5565000:in std_logic;
    clk_logic_5565000:in std_logic;
    m_axis_data_tdata:out std_logic_vector(41 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(24 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_d0050991ffa08d9151315827675f900b;


architecture behavior of xlfir_compiler_d0050991ffa08d9151315827675f900b  is
  component fr_cmplr_v6_3_555df73bebb69ee8
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(47 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(31 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(41 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(41 downto 0);
  s_axis_data_tdata_net(24 downto 0) <= s_axis_data_tdata;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 42,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_11130000,
        clr => '0',
        clk => clk_11130000, 
        o => m_axis_data_tdata
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_11130000,
        clr => '0',
        clk => clk_11130000, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_11130000, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_555df73bebb69ee8_instance : fr_cmplr_v6_3_555df73bebb69ee8
    port map(
      aclk=>clk,
      aclken=>ce_5565000,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_5565000
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_8639b3660dc5b7c78f3b8f56b4679494 is 
  port(
    ce:in std_logic;
    ce_2782500:in std_logic;
    ce_5565000:in std_logic;
    ce_logic_2782500:in std_logic;
    clk:in std_logic;
    clk_2782500:in std_logic;
    clk_5565000:in std_logic;
    clk_logic_2782500:in std_logic;
    m_axis_data_tdata:out std_logic_vector(40 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_8639b3660dc5b7c78f3b8f56b4679494;


architecture behavior of xlfir_compiler_8639b3660dc5b7c78f3b8f56b4679494  is
  component fr_cmplr_v6_3_85eb797d79431254
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(47 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(40 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(40 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 41,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_5565000,
        clr => '0',
        clk => clk_5565000, 
        o => m_axis_data_tdata
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_5565000,
        clr => '0',
        clk => clk_5565000, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_5565000, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_85eb797d79431254_instance : fr_cmplr_v6_3_85eb797d79431254
    port map(
      aclk=>clk,
      aclken=>ce_2782500,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_2782500
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_472d6cb416f02569126e68c627373423 is 
  port(
    ce:in std_logic;
    ce_11130000:in std_logic;
    ce_5565000:in std_logic;
    ce_logic_5565000:in std_logic;
    clk:in std_logic;
    clk_11130000:in std_logic;
    clk_5565000:in std_logic;
    clk_logic_5565000:in std_logic;
    m_axis_data_tdata:out std_logic_vector(42 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(25 downto 0);
    s_axis_data_tready:out std_logic;
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_472d6cb416f02569126e68c627373423;


architecture behavior of xlfir_compiler_472d6cb416f02569126e68c627373423  is
  component fr_cmplr_v6_3_121326a881aa557e
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(47 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(31 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(42 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(42 downto 0);
  s_axis_data_tdata_net(25 downto 0) <= s_axis_data_tdata;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 43,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_11130000,
        clr => '0',
        clk => clk_11130000, 
        o => m_axis_data_tdata
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_11130000,
        clr => '0',
        clk => clk_11130000, 
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_11130000, 
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_121326a881aa557e_instance : fr_cmplr_v6_3_121326a881aa557e
    port map(
      aclk=>clk,
      aclken=>ce_5565000,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_5565000
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_0d0fc5690d is
  port (
    in0 : in std_logic_vector((27 - 1) downto 0);
    in1 : in std_logic_vector((23 - 1) downto 0);
    y : out std_logic_vector((50 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_0d0fc5690d;


architecture behavior of concat_0d0fc5690d is
  signal in0_1_23: unsigned((27 - 1) downto 0);
  signal in1_1_27: unsigned((23 - 1) downto 0);
  signal y_2_1_concat: unsigned((50 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_1d284b35d5 is
  port (
    input_port : in std_logic_vector((50 - 1) downto 0);
    output_port : out std_logic_vector((50 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_1d284b35d5;


architecture behavior of reinterpret_1d284b35d5 is
  signal input_port_1_40: unsigned((50 - 1) downto 0);
  signal output_port_5_5_force: signed((50 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_48a79104f5 is
  port (
    input_port : in std_logic_vector((23 - 1) downto 0);
    output_port : out std_logic_vector((23 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_48a79104f5;


architecture behavior of reinterpret_48a79104f5 is
  signal input_port_1_40: unsigned((23 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_bf9824e821 is
  port (
    input_port : in std_logic_vector((27 - 1) downto 0);
    output_port : out std_logic_vector((27 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_bf9824e821;


architecture behavior of reinterpret_bf9824e821 is
  signal input_port_1_40: signed((27 - 1) downto 0);
  signal output_port_5_5_force: unsigned((27 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity expr_24cbf78c62 is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    c : in std_logic_vector((1 - 1) downto 0);
    d : in std_logic_vector((1 - 1) downto 0);
    dout : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end expr_24cbf78c62;


architecture behavior of expr_24cbf78c62 is
  signal a_1_24: boolean;
  signal b_1_27: boolean;
  signal c_1_30: boolean;
  signal d_1_33: boolean;
  signal bit_7_53: boolean;
  signal bit_7_36: boolean;
  signal fulldout_7_2_bit: boolean;
begin
  a_1_24 <= ((a) = "1");
  b_1_27 <= ((b) = "1");
  c_1_30 <= ((c) = "1");
  d_1_33 <= ((d) = "1");
  bit_7_53 <= ((boolean_to_vector(b_1_27) and boolean_to_vector(a_1_24)) = "1");
  bit_7_36 <= ((boolean_to_vector(c_1_30) and boolean_to_vector(bit_7_53)) = "1");
  fulldout_7_2_bit <= ((boolean_to_vector(d_1_33) and boolean_to_vector(bit_7_36)) = "1");
  dout <= boolean_to_vector(fulldout_7_2_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity expr_375d7bbece is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    c : in std_logic_vector((1 - 1) downto 0);
    dout : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end expr_375d7bbece;


architecture behavior of expr_375d7bbece is
  signal a_1_24: boolean;
  signal b_1_27: boolean;
  signal c_1_30: boolean;
  signal bit_6_36: boolean;
  signal fulldout_6_2_bit: boolean;
begin
  a_1_24 <= ((a) = "1");
  b_1_27 <= ((b) = "1");
  c_1_30 <= ((c) = "1");
  bit_6_36 <= ((boolean_to_vector(b_1_27) and boolean_to_vector(a_1_24)) = "1");
  fulldout_6_2_bit <= ((boolean_to_vector(c_1_30) and boolean_to_vector(bit_6_36)) = "1");
  dout <= boolean_to_vector(fulldout_6_2_bit);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.conv_pkg.all;
entity xlfifogen is
  generic (
    core_name0: string := "";
    data_width: integer := -1;
    data_count_width: integer := -1;
    percent_full_width: integer := -1;
    has_ae : integer := 0;
    has_af : integer := 0
  );
  port (
    din: in std_logic_vector(data_width - 1 downto 0);
    we: in std_logic;
    we_ce: in std_logic;
    re: in std_logic;
    re_ce: in std_logic;
    rst: in std_logic;
    en: in std_logic;
    ce: in std_logic;
    clk: in std_logic;
    empty: out std_logic;
    full: out std_logic;
    percent_full: out std_logic_vector(percent_full_width - 1 downto 0);
    dcount: out std_logic_vector(data_count_width - 1 downto 0);
    ae: out std_logic;
    af: out std_logic;
    dout: out std_logic_vector(data_width - 1 downto 0)
  );
end xlfifogen ;
architecture behavior of xlfifogen is
  component fifo_fg84_26bc5f646d342e7f
    port (
      clk: in std_logic;
      din: in std_logic_vector(data_width - 1 downto 0);
      wr_en: in std_logic;
      rd_en: in std_logic;
      dout: out std_logic_vector(data_width - 1 downto 0);
      full: out std_logic;
      empty: out std_logic
    );
  end component;
  attribute syn_black_box of fifo_fg84_26bc5f646d342e7f:
    component is true;
  attribute fpga_dont_touch of fifo_fg84_26bc5f646d342e7f:
    component is "true";
  attribute box_type of fifo_fg84_26bc5f646d342e7f:
    component  is "black_box";
  signal rd_en: std_logic;
  signal wr_en: std_logic;
  signal srst: std_logic;
  signal core_full: std_logic;
  signal core_dcount: std_logic_vector(data_count_width - 1 downto 0);
begin
  comp0: if ((core_name0 = "fifo_fg84_26bc5f646d342e7f")) generate
    core_instance0: fifo_fg84_26bc5f646d342e7f
      port map (
        clk => clk,
        din => din,
        wr_en => wr_en,
        rd_en => rd_en,
        dout => dout,
        full => core_full,
        empty => empty
      );
  end generate;

  modify_count: process(core_full, core_dcount) is
  begin
    if core_full = '1' then
      percent_full <= (others => '1');
    else
      percent_full <= core_dcount(data_count_width-1 downto data_count_width-percent_full_width);
    end if;
  end process modify_count;

  rd_en <= re and en and re_ce;
  wr_en <= we and en and we_ce;
  full <= core_full;
  srst <= rst and ce;
  dcount <= core_dcount;

  terminate_core_ae: if has_ae /= 1 generate
  begin
    ae <= '0';
  end generate terminate_core_ae;
  terminate_core_af: if has_af /= 1 generate
  begin
    af <= '0';
  end generate terminate_core_af;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_fractional:out std_logic_vector(22 downto 0);
    m_axis_dout_tdata_quotient:out std_logic_vector(26 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_dividend_tdata_dividend:in std_logic_vector(26 downto 0);
    s_axis_dividend_tready:out std_logic;
    s_axis_dividend_tvalid:in std_logic;
    s_axis_divisor_tdata_divisor:in std_logic_vector(26 downto 0);
    s_axis_divisor_tready:out std_logic;
    s_axis_divisor_tvalid:in std_logic
  );
end xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7;


architecture behavior of xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7  is
  component dv_gn_v4_0_5ce7b020ea0b7ee9
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(79 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_dividend_tdata:in std_logic_vector(31 downto 0);
      s_axis_dividend_tready:out std_logic;
      s_axis_dividend_tvalid:in std_logic;
      s_axis_divisor_tdata:in std_logic_vector(31 downto 0);
      s_axis_divisor_tready:out std_logic;
      s_axis_divisor_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(79 downto 0) := (others=>'0');
signal m_axis_dout_tdata_quotient_net: std_logic_vector(26 downto 0) := (others=>'0');
signal m_axis_dout_tdata_shift_out_net: std_logic_vector(49 downto 0) := (others=>'0');
signal m_axis_dout_tdata_fractional_net: std_logic_vector(45 downto 0) := (others=>'0');
signal s_axis_dividend_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal s_axis_divisor_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_quotient_net <= m_axis_dout_tdata_net(72 downto 46);
  m_axis_dout_tdata_fractional_net <= m_axis_dout_tdata_net(45 downto 0);
  s_axis_dividend_tdata_net(26 downto 0) <= s_axis_dividend_tdata_dividend;
  s_axis_divisor_tdata_net(26 downto 0) <= s_axis_divisor_tdata_divisor;
  m_axis_dout_tdata_quotient <= m_axis_dout_tdata_shift_out_net(49 downto 23);
m_axis_dout_tdata_fractional <= m_axis_dout_tdata_shift_out_net(22 downto 0);
m_axis_dout_tdata_shift_out_net <= shift_division_result(m_axis_dout_tdata_quotient_net, m_axis_dout_tdata_fractional_net, 23, 0, 1);
  dv_gn_v4_0_5ce7b020ea0b7ee9_instance : dv_gn_v4_0_5ce7b020ea0b7ee9
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_dividend_tdata=>s_axis_dividend_tdata_net,
      s_axis_dividend_tready=>s_axis_dividend_tready,
      s_axis_dividend_tvalid=>s_axis_dividend_tvalid,
      s_axis_divisor_tdata=>s_axis_divisor_tdata_net,
      s_axis_divisor_tready=>s_axis_divisor_tready,
      s_axis_divisor_tvalid=>s_axis_divisor_tvalid
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6505656e93 is
  port (
    a : in std_logic_vector((27 - 1) downto 0);
    b : in std_logic_vector((27 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6505656e93;


architecture behavior of relational_6505656e93 is
  signal a_1_31: signed((27 - 1) downto 0);
  signal b_1_34: signed((27 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_signed(a);
  b_1_34 <= std_logic_vector_to_signed(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub;
architecture behavior of xladdsub is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_239e4f614ba09ab1
    port (
          a: in std_logic_vector(26 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(26 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_239e4f614ba09ab1:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_239e4f614ba09ab1:
    component is "true";
  attribute box_type of addsb_11_0_239e4f614ba09ab1:
    component  is "black_box";
  component addsb_11_0_1482f9e8df81448a
    port (
          a: in std_logic_vector(27 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(27 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_1482f9e8df81448a:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_1482f9e8df81448a:
    component is "true";
  attribute box_type of addsb_11_0_1482f9e8df81448a:
    component  is "black_box";
  component addsb_11_0_2f1626aeedb3c308
    port (
          a: in std_logic_vector(27 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(27 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_2f1626aeedb3c308:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_2f1626aeedb3c308:
    component is "true";
  attribute box_type of addsb_11_0_2f1626aeedb3c308:
    component  is "black_box";
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_239e4f614ba09ab1")) generate
    core_instance0: addsb_11_0_239e4f614ba09ab1
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp1: if ((core_name0 = "addsb_11_0_1482f9e8df81448a")) generate
    core_instance1: addsb_11_0_1482f9e8df81448a
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_2f1626aeedb3c308")) generate
    core_instance2: addsb_11_0_2f1626aeedb3c308
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xldds_compiler_b7bbc719459e4bb4074716a9175f7d86 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_data_tdata_cosine:out std_logic_vector(23 downto 0);
    m_axis_data_tdata_sine:out std_logic_vector(23 downto 0);
    m_axis_data_tready:in std_logic;
    m_axis_data_tvalid:out std_logic
  );
end xldds_compiler_b7bbc719459e4bb4074716a9175f7d86;


architecture behavior of xldds_compiler_b7bbc719459e4bb4074716a9175f7d86  is
  component dds_cmplr_v5_0_61b575ede3cdcc97
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_data_tdata:out std_logic_vector(47 downto 0);
      m_axis_data_tready:in std_logic;
      m_axis_data_tvalid:out std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_sine <= m_axis_data_tdata_net(47 downto 24);
  m_axis_data_tdata_cosine <= m_axis_data_tdata_net(23 downto 0);
  dds_cmplr_v5_0_61b575ede3cdcc97_instance : dds_cmplr_v5_0_61b575ede3cdcc97
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tready=>m_axis_data_tready,
      m_axis_data_tvalid=>m_axis_data_tvalid
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xldsamp is
  generic (
    d_width: integer := 12;
    d_bin_pt: integer := 0;
    d_arith: integer := xlUnsigned;
    q_width: integer := 12;
    q_bin_pt: integer := 0;
    q_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    ds_ratio: integer := 2;
    phase: integer := 0;
    latency: integer := 1
  );
  port (
    d: in std_logic_vector(d_width - 1 downto 0);
    src_clk: in std_logic;
    src_ce: in std_logic;
    src_clr: in std_logic;
    dest_clk: in std_logic;
    dest_ce: in std_logic;
    dest_clr: in std_logic;
    en: in std_logic_vector(en_width - 1 downto 0);
    q: out std_logic_vector(q_width - 1 downto 0)
  );
end xldsamp;
architecture struct of xldsamp is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component fdse
    port (
      q: out   std_ulogic;
      d: in    std_ulogic;
      c: in    std_ulogic;
      s: in    std_ulogic;
      ce: in    std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  signal adjusted_dest_ce: std_logic;
  signal adjusted_dest_ce_w_en: std_logic;
  signal dest_ce_w_en: std_logic;
  signal smpld_d: std_logic_vector(d_width-1 downto 0);
begin
  adjusted_ce_needed: if ((latency = 0) or (phase /= (ds_ratio - 1))) generate
    dest_ce_reg: fdse
      port map (
        q => adjusted_dest_ce,
        d => dest_ce,
        c => src_clk,
        s => src_clr,
        ce => src_ce
      );
  end generate;
  latency_eq_0: if (latency = 0) generate
    shutter_d_reg: synth_reg
      generic map (
        width => d_width,
        latency => 1
      )
      port map (
        i => d,
        ce => adjusted_dest_ce,
        clr => src_clr,
        clk => src_clk,
        o => smpld_d
      );
    shutter_mux: process (adjusted_dest_ce, d, smpld_d)
    begin
      if adjusted_dest_ce = '0' then
        q <= smpld_d;
      else
        q <= d;
      end if;
    end process;
  end generate;
  latency_gt_0: if (latency > 0) generate
    dbl_reg_test: if (phase /= (ds_ratio-1)) generate
        smpl_d_reg: synth_reg
          generic map (
            width => d_width,
            latency => 1
          )
          port map (
            i => d,
            ce => adjusted_dest_ce_w_en,
            clr => src_clr,
            clk => src_clk,
            o => smpld_d
          );
    end generate;
    sngl_reg_test: if (phase = (ds_ratio -1)) generate
      smpld_d <= d;
    end generate;
    latency_pipe: synth_reg
      generic map (
        width => d_width,
        latency => latency
      )
      port map (
        i => smpld_d,
        ce => dest_ce_w_en,
        clr => src_clr,
        clk => dest_clk,
        o => q
      );
  end generate;
  dest_ce_w_en <= dest_ce and en(0);
  adjusted_dest_ce_w_en <= adjusted_dest_ce and en(0);
end architecture struct;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_fofb/cic_fofb"

entity cic_fofb_entity_c0b771be35 is
  port (
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    i_in: in std_logic_vector(23 downto 0); 
    q_in: in std_logic_vector(23 downto 0); 
    i_out: out std_logic_vector(24 downto 0); 
    i_valid: out std_logic; 
    q_out: out std_logic_vector(24 downto 0)
  );
end cic_fofb_entity_c0b771be35;

architecture structural of cic_fofb_entity_c0b771be35 is
  signal ce_1113_sg_x0: std_logic;
  signal ce_1_sg_x0: std_logic;
  signal ce_logic_1_sg_x0: std_logic;
  signal cic_fofb_i_m_axis_data_tdata_data_net: std_logic_vector(24 downto 0);
  signal cic_fofb_i_m_axis_data_tvalid_net_x0: std_logic;
  signal cic_fofb_q_m_axis_data_tdata_data_net: std_logic_vector(24 downto 0);
  signal clk_1113_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal delay6_q_net_x0: std_logic_vector(23 downto 0);
  signal delay7_q_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  ce_1113_sg_x0 <= ce_1113;
  ce_logic_1_sg_x0 <= ce_logic_1;
  clk_1_sg_x0 <= clk_1;
  clk_1113_sg_x0 <= clk_1113;
  delay7_q_net_x0 <= i_in;
  delay6_q_net_x0 <= q_in;
  i_out <= reinterpret1_output_port_net_x0;
  i_valid <= cic_fofb_i_m_axis_data_tvalid_net_x0;
  q_out <= reinterpret_output_port_net_x0;

  cic_fofb_i: entity work.xlcic_compiler_bb7d6f586f04abec4d028ced88abc8ae
    port map (
      ce => ce_1_sg_x0,
      ce_1113 => ce_1113_sg_x0,
      ce_logic_1 => ce_logic_1_sg_x0,
      clk => clk_1_sg_x0,
      clk_1113 => clk_1113_sg_x0,
      clk_logic_1 => clk_1_sg_x0,
      s_axis_data_tdata_data => delay7_q_net_x0,
      m_axis_data_tdata_data => cic_fofb_i_m_axis_data_tdata_data_net,
      m_axis_data_tvalid => cic_fofb_i_m_axis_data_tvalid_net_x0
    );

  cic_fofb_q: entity work.xlcic_compiler_bb7d6f586f04abec4d028ced88abc8ae
    port map (
      ce => ce_1_sg_x0,
      ce_1113 => ce_1113_sg_x0,
      ce_logic_1 => ce_logic_1_sg_x0,
      clk => clk_1_sg_x0,
      clk_1113 => clk_1113_sg_x0,
      clk_logic_1 => clk_1_sg_x0,
      s_axis_data_tdata_data => delay6_q_net_x0,
      m_axis_data_tdata_data => cic_fofb_q_m_axis_data_tdata_data_net
    );

  reinterpret: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_fofb_q_m_axis_data_tdata_data_net,
      output_port => reinterpret_output_port_net_x0
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_fofb_i_m_axis_data_tdata_data_net,
      output_port => reinterpret1_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_fofb"

entity channel0_fofb_entity_3577a252e5 is
  port (
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    mix_i_in: in std_logic_vector(23 downto 0); 
    mix_q_in: in std_logic_vector(23 downto 0); 
    amp_f: out std_logic_vector(24 downto 0); 
    cic_fofb_i_fpga_out: out std_logic_vector(24 downto 0); 
    cic_fofb_q_fpga_out: out std_logic_vector(24 downto 0); 
    valid_f: out std_logic
  );
end channel0_fofb_entity_3577a252e5;

architecture structural of channel0_fofb_entity_3577a252e5 is
  signal ce_1113_sg_x1: std_logic;
  signal ce_1_sg_x1: std_logic;
  signal ce_logic_1_sg_x1: std_logic;
  signal cic_fofb_i_m_axis_data_tvalid_net_x0: std_logic;
  signal clk_1113_sg_x1: std_logic;
  signal clk_1_sg_x1: std_logic;
  signal delay6_q_net_x1: std_logic_vector(23 downto 0);
  signal delay7_q_net_x1: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(24 downto 0);
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register5_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal reinterpret1_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x1: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x1 <= ce_1;
  ce_1113_sg_x1 <= ce_1113;
  ce_logic_1_sg_x1 <= ce_logic_1;
  clk_1_sg_x1 <= clk_1;
  clk_1113_sg_x1 <= clk_1113;
  delay7_q_net_x1 <= mix_i_in;
  delay6_q_net_x1 <= mix_q_in;
  amp_f <= register5_q_net_x0;
  cic_fofb_i_fpga_out <= reinterpret1_output_port_net_x1;
  cic_fofb_q_fpga_out <= reinterpret_output_port_net_x1;
  valid_f <= register6_q_net_x0;

  cic_fofb_c0b771be35: entity work.cic_fofb_entity_c0b771be35
    port map (
      ce_1 => ce_1_sg_x1,
      ce_1113 => ce_1113_sg_x1,
      ce_logic_1 => ce_logic_1_sg_x1,
      clk_1 => clk_1_sg_x1,
      clk_1113 => clk_1113_sg_x1,
      i_in => delay7_q_net_x1,
      q_in => delay6_q_net_x1,
      i_out => reinterpret1_output_port_net_x1,
      i_valid => cic_fofb_i_m_axis_data_tvalid_net_x0,
      q_out => reinterpret_output_port_net_x1
    );

  rect2pol: entity work.xlcordic_c062cc3a2d77ede2032de397150e15cd
    port map (
      ce => ce_1113_sg_x1,
      clk => clk_1113_sg_x1,
      s_axis_cartesian_tdata_imag => reinterpret_output_port_net_x1,
      s_axis_cartesian_tdata_real => reinterpret1_output_port_net_x1,
      s_axis_cartesian_tvalid => cic_fofb_i_m_axis_data_tvalid_net_x0,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x1,
      clk => clk_1113_sg_x1,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1113_sg_x1,
      clk => clk_1113_sg_x1,
      d(0) => rect2pol_m_axis_dout_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt/DDC/DataReg_En"

entity datareg_en_entity_3ccf612162 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(23 downto 0); 
    en: in std_logic; 
    dout: out std_logic_vector(23 downto 0)
  );
end datareg_en_entity_3ccf612162;

architecture structural of datareg_en_entity_3ccf612162 is
  signal bpf_fpga_m_axis_data_tvalid_net_x0: std_logic;
  signal ce_1_sg_x2: std_logic;
  signal clk_1_sg_x2: std_logic;
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x0: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x2 <= ce_1;
  clk_1_sg_x2 <= clk_1;
  convert_dout_net_x0 <= din;
  bpf_fpga_m_axis_data_tvalid_net_x0 <= en;
  dout <= register_q_net_x0;

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x2,
      clk => clk_1_sg_x2,
      d => convert_dout_net_x0,
      en(0) => bpf_fpga_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt/DDC/Mixer/DataReg_En"

entity datareg_en_entity_c073dad362 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    din: in std_logic_vector(23 downto 0); 
    en: in std_logic; 
    dout: out std_logic_vector(23 downto 0); 
    valid: out std_logic
  );
end datareg_en_entity_c073dad362;

architecture structural of datareg_en_entity_c073dad362 is
  signal ce_1_sg_x3: std_logic;
  signal clk_1_sg_x3: std_logic;
  signal constant1_op_net_x0: std_logic;
  signal constant2_op_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x3 <= ce_1;
  clk_1_sg_x3 <= clk_1;
  constant2_op_net_x0 <= din;
  constant1_op_net_x0 <= en;
  dout <= register_q_net_x0;
  valid <= register1_q_net_x0;

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      d(0) => constant1_op_net_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      d => constant2_op_net_x0,
      en(0) => constant1_op_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt/DDC/Mixer"

entity mixer_entity_9216a510d2 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    dds_cosine: in std_logic_vector(23 downto 0); 
    dds_msine: in std_logic_vector(23 downto 0); 
    dds_valid: in std_logic; 
    din_i: in std_logic_vector(23 downto 0); 
    din_q: in std_logic_vector(23 downto 0); 
    en: in std_logic; 
    i: out std_logic_vector(23 downto 0); 
    q: out std_logic_vector(23 downto 0)
  );
end mixer_entity_9216a510d2;

architecture structural of mixer_entity_9216a510d2 is
  signal a_i: std_logic_vector(23 downto 0);
  signal a_r: std_logic_vector(23 downto 0);
  signal b_i: std_logic_vector(23 downto 0);
  signal b_r: std_logic_vector(23 downto 0);
  signal ce_1_sg_x5: std_logic;
  signal clk_1_sg_x5: std_logic;
  signal complexmult_m_axis_dout_tdata_imag_net: std_logic_vector(23 downto 0);
  signal complexmult_m_axis_dout_tdata_real_net: std_logic_vector(23 downto 0);
  signal complexmult_m_axis_dout_tvalid_net: std_logic;
  signal constant1_op_net_x2: std_logic;
  signal constant2_op_net_x1: std_logic_vector(23 downto 0);
  signal convert1_dout_net: std_logic_vector(23 downto 0);
  signal convert2_dout_net: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x0: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x0: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x0: std_logic;
  signal delay6_q_net_x2: std_logic_vector(23 downto 0);
  signal delay7_q_net_x2: std_logic_vector(23 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x2: std_logic_vector(23 downto 0);
  signal register_q_net_x3: std_logic_vector(23 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x5 <= ce_1;
  clk_1_sg_x5 <= clk_1;
  dds_m_axis_data_tdata_cosine_net_x0 <= dds_cosine;
  dds_m_axis_data_tdata_sine_net_x0 <= dds_msine;
  dds_m_axis_data_tvalid_net_x0 <= dds_valid;
  register_q_net_x3 <= din_i;
  constant2_op_net_x1 <= din_q;
  constant1_op_net_x2 <= en;
  i <= delay7_q_net_x2;
  q <= delay6_q_net_x2;

  complexmult: entity work.xlcomplex_multiplier_a3a52a268f0fdc1111e428e7f4c7c82c
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      s_axis_a_tdata_imag => a_i,
      s_axis_a_tdata_real => a_r,
      s_axis_a_tvalid => dds_m_axis_data_tvalid_net_x0,
      s_axis_b_tdata_imag => b_i,
      s_axis_b_tdata_real => b_r,
      s_axis_b_tvalid => register1_q_net_x0,
      m_axis_dout_tdata_imag => complexmult_m_axis_dout_tdata_imag_net,
      m_axis_dout_tdata_real => complexmult_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => complexmult_m_axis_dout_tvalid_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 19,
      din_width => 24,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      clr => '0',
      din => reinterpret1_output_port_net,
      en => "1",
      dout => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 19,
      din_width => 24,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert2_dout_net
    );

  datareg_en1_02ef0305a4: entity work.datareg_en_entity_3ccf612162
    port map (
      ce_1 => ce_1_sg_x5,
      clk_1 => clk_1_sg_x5,
      din => register_q_net_x3,
      en => constant1_op_net_x2,
      dout => register_q_net_x2
    );

  datareg_en_c073dad362: entity work.datareg_en_entity_c073dad362
    port map (
      ce_1 => ce_1_sg_x5,
      clk_1 => clk_1_sg_x5,
      din => constant2_op_net_x1,
      en => constant1_op_net_x2,
      dout => register_q_net_x0,
      valid => register1_q_net_x0
    );

  delay: entity work.delay_961b43f67a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => register_q_net_x0,
      q => b_i
    );

  delay1: entity work.delay_961b43f67a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => register_q_net_x2,
      q => b_r
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      d => dds_m_axis_data_tdata_sine_net_x0,
      en => dds_m_axis_data_tvalid_net_x0,
      rst => '1',
      q => a_i
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      d => dds_m_axis_data_tdata_cosine_net_x0,
      en => dds_m_axis_data_tvalid_net_x0,
      rst => '1',
      q => a_r
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      d => convert2_dout_net,
      en => complexmult_m_axis_dout_tvalid_net,
      rst => '1',
      q => delay6_q_net_x2
    );

  delay7: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      d => convert1_dout_net,
      en => complexmult_m_axis_dout_tvalid_net,
      rst => '1',
      q => delay7_q_net_x2
    );

  reinterpret: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => complexmult_m_axis_dout_tdata_imag_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => complexmult_m_axis_dout_tdata_real_net,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt/DDC"

entity ddc_entity_fbec30928b is
  port (
    adc_in: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    dds_cosine_in: in std_logic_vector(23 downto 0); 
    dds_msine_in: in std_logic_vector(23 downto 0); 
    dds_valid_in: in std_logic; 
    bpf_out: out std_logic_vector(23 downto 0); 
    mix_i_out: out std_logic_vector(23 downto 0); 
    mix_q_out: out std_logic_vector(23 downto 0)
  );
end ddc_entity_fbec30928b;

architecture structural of ddc_entity_fbec30928b is
  signal adc_ch0_i_net_x0: std_logic_vector(15 downto 0);
  signal bpf_fpga_m_axis_data_tdata_net: std_logic_vector(33 downto 0);
  signal bpf_fpga_m_axis_data_tvalid_net_x0: std_logic;
  signal ce_1_sg_x6: std_logic;
  signal ce_logic_1_sg_x2: std_logic;
  signal clk_1_sg_x6: std_logic;
  signal constant1_op_net_x2: std_logic;
  signal constant2_op_net_x1: std_logic_vector(23 downto 0);
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x1: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x1: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x1: std_logic;
  signal delay6_q_net_x3: std_logic_vector(23 downto 0);
  signal delay7_q_net_x3: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(15 downto 0);
  signal register_q_net_x4: std_logic_vector(23 downto 0);

begin
  adc_ch0_i_net_x0 <= adc_in;
  ce_1_sg_x6 <= ce_1;
  ce_logic_1_sg_x2 <= ce_logic_1;
  clk_1_sg_x6 <= clk_1;
  dds_m_axis_data_tdata_cosine_net_x1 <= dds_cosine_in;
  dds_m_axis_data_tdata_sine_net_x1 <= dds_msine_in;
  dds_m_axis_data_tvalid_net_x1 <= dds_valid_in;
  bpf_out <= register_q_net_x4;
  mix_i_out <= delay7_q_net_x3;
  mix_q_out <= delay6_q_net_x3;

  bpf_fpga: entity work.xlfir_compiler_db690cb1dac026c47ff98d5afcede74f
    port map (
      ce => ce_1_sg_x6,
      ce_logic_1 => ce_logic_1_sg_x2,
      clk => clk_1_sg_x6,
      clk_logic_1 => clk_1_sg_x6,
      s_axis_data_tdata => register_q_net,
      src_ce => ce_1_sg_x6,
      src_clk => clk_1_sg_x6,
      m_axis_data_tdata => bpf_fpga_m_axis_data_tdata_net,
      m_axis_data_tvalid => bpf_fpga_m_axis_data_tvalid_net_x0
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net_x2
    );

  constant2: entity work.constant_f394f3309c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net_x1
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 32,
      din_width => 34,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      din => bpf_fpga_m_axis_data_tdata_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  datareg_en_3ccf612162: entity work.datareg_en_entity_3ccf612162
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      din => convert_dout_net_x0,
      en => bpf_fpga_m_axis_data_tvalid_net_x0,
      dout => register_q_net_x4
    );

  mixer_9216a510d2: entity work.mixer_entity_9216a510d2
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      dds_cosine => dds_m_axis_data_tdata_cosine_net_x1,
      dds_msine => dds_m_axis_data_tdata_sine_net_x1,
      dds_valid => dds_m_axis_data_tvalid_net_x1,
      din_i => register_q_net_x4,
      din_q => constant2_op_net_x1,
      en => constant1_op_net_x2,
      i => delay7_q_net_x3,
      q => delay6_q_net_x3
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      d => adc_ch0_i_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt/decim35"

entity decim35_entity_3519cdb9ab is
  port (
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    i_in: in std_logic_vector(23 downto 0); 
    q_in: in std_logic_vector(23 downto 0); 
    i_out: out std_logic_vector(24 downto 0); 
    q_out: out std_logic_vector(24 downto 0); 
    valid_out: out std_logic
  );
end decim35_entity_3519cdb9ab;

architecture structural of decim35_entity_3519cdb9ab is
  signal ce_1_sg_x7: std_logic;
  signal ce_35_sg_x0: std_logic;
  signal ce_logic_1_sg_x3: std_logic;
  signal clk_1_sg_x7: std_logic;
  signal clk_35_sg_x0: std_logic;
  signal convert1_dout_net_x0: std_logic_vector(24 downto 0);
  signal convert2_dout_net_x0: std_logic_vector(24 downto 0);
  signal delay6_q_net_x4: std_logic_vector(23 downto 0);
  signal delay7_q_net_x4: std_logic_vector(23 downto 0);
  signal fir_compiler_6_2_m_axis_data_tdata_path0_net: std_logic_vector(44 downto 0);
  signal fir_compiler_6_2_m_axis_data_tdata_path1_net: std_logic_vector(44 downto 0);
  signal fir_compiler_6_2_m_axis_data_tvalid_net_x0: std_logic;
  signal reinterpret1_output_port_net: std_logic_vector(44 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(44 downto 0);

begin
  ce_1_sg_x7 <= ce_1;
  ce_35_sg_x0 <= ce_35;
  ce_logic_1_sg_x3 <= ce_logic_1;
  clk_1_sg_x7 <= clk_1;
  clk_35_sg_x0 <= clk_35;
  delay7_q_net_x4 <= i_in;
  delay6_q_net_x4 <= q_in;
  i_out <= convert2_dout_net_x0;
  q_out <= convert1_dout_net_x0;
  valid_out <= fir_compiler_6_2_m_axis_data_tvalid_net_x0;

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 42,
      din_width => 45,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert1_dout_net_x0
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 42,
      din_width => 45,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      clr => '0',
      din => reinterpret1_output_port_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  fir_compiler_6_2: entity work.xlfir_compiler_6d27a36d02c91c0ddc9d14d956c5aca1
    port map (
      ce => ce_1_sg_x7,
      ce_35 => ce_35_sg_x0,
      ce_logic_1 => ce_logic_1_sg_x3,
      clk => clk_1_sg_x7,
      clk_35 => clk_35_sg_x0,
      clk_logic_1 => clk_1_sg_x7,
      s_axis_data_tdata_path0 => delay7_q_net_x4,
      s_axis_data_tdata_path1 => delay6_q_net_x4,
      src_ce => ce_1_sg_x7,
      src_clk => clk_1_sg_x7,
      m_axis_data_tdata_path0 => fir_compiler_6_2_m_axis_data_tdata_path0_net,
      m_axis_data_tdata_path1 => fir_compiler_6_2_m_axis_data_tdata_path1_net,
      m_axis_data_tvalid => fir_compiler_6_2_m_axis_data_tvalid_net_x0
    );

  reinterpret: entity work.reinterpret_82c3c799ff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => fir_compiler_6_2_m_axis_data_tdata_path1_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_82c3c799ff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => fir_compiler_6_2_m_axis_data_tdata_path0_net,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel0_tbt"

entity channel0_tbt_entity_b3ebb9eccb is
  port (
    adc_ch0_i: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    dds_cosine_in: in std_logic_vector(23 downto 0); 
    dds_msine_in: in std_logic_vector(23 downto 0); 
    dds_valid_in: in std_logic; 
    amp_f: out std_logic_vector(24 downto 0); 
    bpf_adc_fpga_out: out std_logic_vector(23 downto 0); 
    decim_35_i_fpga_out: out std_logic_vector(24 downto 0); 
    decim_35_q_fpga_out: out std_logic_vector(24 downto 0); 
    mix_i: out std_logic_vector(23 downto 0); 
    mix_q: out std_logic_vector(23 downto 0); 
    valid_f: out std_logic
  );
end channel0_tbt_entity_b3ebb9eccb;

architecture structural of channel0_tbt_entity_b3ebb9eccb is
  signal adc_ch0_i_net_x1: std_logic_vector(15 downto 0);
  signal ce_1_sg_x8: std_logic;
  signal ce_35_sg_x1: std_logic;
  signal ce_logic_1_sg_x4: std_logic;
  signal clk_1_sg_x8: std_logic;
  signal clk_35_sg_x1: std_logic;
  signal convert1_dout_net_x1: std_logic_vector(24 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(24 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x2: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x2: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x2: std_logic;
  signal delay6_q_net_x5: std_logic_vector(23 downto 0);
  signal delay7_q_net_x5: std_logic_vector(23 downto 0);
  signal fir_compiler_6_2_m_axis_data_tvalid_net_x0: std_logic;
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(24 downto 0);
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register5_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal register_q_net_x5: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);

begin
  adc_ch0_i_net_x1 <= adc_ch0_i;
  ce_1_sg_x8 <= ce_1;
  ce_35_sg_x1 <= ce_35;
  ce_logic_1_sg_x4 <= ce_logic_1;
  clk_1_sg_x8 <= clk_1;
  clk_35_sg_x1 <= clk_35;
  dds_m_axis_data_tdata_cosine_net_x2 <= dds_cosine_in;
  dds_m_axis_data_tdata_sine_net_x2 <= dds_msine_in;
  dds_m_axis_data_tvalid_net_x2 <= dds_valid_in;
  amp_f <= register5_q_net_x0;
  bpf_adc_fpga_out <= register_q_net_x5;
  decim_35_i_fpga_out <= convert2_dout_net_x1;
  decim_35_q_fpga_out <= convert1_dout_net_x1;
  mix_i <= delay7_q_net_x5;
  mix_q <= delay6_q_net_x5;
  valid_f <= register6_q_net_x0;

  ddc_fbec30928b: entity work.ddc_entity_fbec30928b
    port map (
      adc_in => adc_ch0_i_net_x1,
      ce_1 => ce_1_sg_x8,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x8,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x2,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x2,
      dds_valid_in => dds_m_axis_data_tvalid_net_x2,
      bpf_out => register_q_net_x5,
      mix_i_out => delay7_q_net_x5,
      mix_q_out => delay6_q_net_x5
    );

  decim35_3519cdb9ab: entity work.decim35_entity_3519cdb9ab
    port map (
      ce_1 => ce_1_sg_x8,
      ce_35 => ce_35_sg_x1,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x8,
      clk_35 => clk_35_sg_x1,
      i_in => delay7_q_net_x5,
      q_in => delay6_q_net_x5,
      i_out => convert2_dout_net_x1,
      q_out => convert1_dout_net_x1,
      valid_out => fir_compiler_6_2_m_axis_data_tvalid_net_x0
    );

  rect2pol: entity work.xlcordic_c062cc3a2d77ede2032de397150e15cd
    port map (
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      s_axis_cartesian_tdata_imag => convert1_dout_net_x1,
      s_axis_cartesian_tdata_real => convert2_dout_net_x1,
      s_axis_cartesian_tvalid => fir_compiler_6_2_m_axis_data_tvalid_net_x0,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      d(0) => rect2pol_m_axis_dout_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel1_tbt"

entity channel1_tbt_entity_8d468f1125 is
  port (
    adc_ch1_i: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    dds_cosine_in: in std_logic_vector(23 downto 0); 
    dds_msine_in: in std_logic_vector(23 downto 0); 
    dds_valid_in: in std_logic; 
    amp_f: out std_logic_vector(24 downto 0); 
    bpf_adc_fpga_out: out std_logic_vector(23 downto 0); 
    decim_35_i_fpga_out: out std_logic_vector(24 downto 0); 
    decim_35_q_fpga_out: out std_logic_vector(24 downto 0); 
    mix_i: out std_logic_vector(23 downto 0); 
    mix_q: out std_logic_vector(23 downto 0); 
    valid_f: out std_logic
  );
end channel1_tbt_entity_8d468f1125;

architecture structural of channel1_tbt_entity_8d468f1125 is
  signal adc_ch1_i_net_x1: std_logic_vector(15 downto 0);
  signal ce_1_sg_x17: std_logic;
  signal ce_35_sg_x3: std_logic;
  signal ce_logic_1_sg_x9: std_logic;
  signal clk_1_sg_x17: std_logic;
  signal clk_35_sg_x3: std_logic;
  signal convert1_dout_net_x1: std_logic_vector(24 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(24 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x5: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x5: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x5: std_logic;
  signal delay6_q_net_x5: std_logic_vector(23 downto 0);
  signal delay7_q_net_x5: std_logic_vector(23 downto 0);
  signal fir_compiler_6_2_m_axis_data_tvalid_net_x0: std_logic;
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(24 downto 0);
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register5_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal register_q_net_x5: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);

begin
  adc_ch1_i_net_x1 <= adc_ch1_i;
  ce_1_sg_x17 <= ce_1;
  ce_35_sg_x3 <= ce_35;
  ce_logic_1_sg_x9 <= ce_logic_1;
  clk_1_sg_x17 <= clk_1;
  clk_35_sg_x3 <= clk_35;
  dds_m_axis_data_tdata_cosine_net_x5 <= dds_cosine_in;
  dds_m_axis_data_tdata_sine_net_x5 <= dds_msine_in;
  dds_m_axis_data_tvalid_net_x5 <= dds_valid_in;
  amp_f <= register5_q_net_x0;
  bpf_adc_fpga_out <= register_q_net_x5;
  decim_35_i_fpga_out <= convert2_dout_net_x1;
  decim_35_q_fpga_out <= convert1_dout_net_x1;
  mix_i <= delay7_q_net_x5;
  mix_q <= delay6_q_net_x5;
  valid_f <= register6_q_net_x0;

  ddc_6518856b7b: entity work.ddc_entity_fbec30928b
    port map (
      adc_in => adc_ch1_i_net_x1,
      ce_1 => ce_1_sg_x17,
      ce_logic_1 => ce_logic_1_sg_x9,
      clk_1 => clk_1_sg_x17,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x5,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x5,
      dds_valid_in => dds_m_axis_data_tvalid_net_x5,
      bpf_out => register_q_net_x5,
      mix_i_out => delay7_q_net_x5,
      mix_q_out => delay6_q_net_x5
    );

  decim35_aa72de60bf: entity work.decim35_entity_3519cdb9ab
    port map (
      ce_1 => ce_1_sg_x17,
      ce_35 => ce_35_sg_x3,
      ce_logic_1 => ce_logic_1_sg_x9,
      clk_1 => clk_1_sg_x17,
      clk_35 => clk_35_sg_x3,
      i_in => delay7_q_net_x5,
      q_in => delay6_q_net_x5,
      i_out => convert2_dout_net_x1,
      q_out => convert1_dout_net_x1,
      valid_out => fir_compiler_6_2_m_axis_data_tvalid_net_x0
    );

  rect2pol: entity work.xlcordic_c062cc3a2d77ede2032de397150e15cd
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      s_axis_cartesian_tdata_imag => convert1_dout_net_x1,
      s_axis_cartesian_tdata_real => convert2_dout_net_x1,
      s_axis_cartesian_tvalid => fir_compiler_6_2_m_axis_data_tvalid_net_x0,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      d(0) => rect2pol_m_axis_dout_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel2_tbt"

entity channel2_tbt_entity_c5e2abdcfa is
  port (
    adc_ch2_i: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    dds_cosine_in: in std_logic_vector(23 downto 0); 
    dds_msine_in: in std_logic_vector(23 downto 0); 
    dds_valid_in: in std_logic; 
    amp_f: out std_logic_vector(24 downto 0); 
    bpf_adc_fpga_out: out std_logic_vector(23 downto 0); 
    decim_35_i_fpga_out: out std_logic_vector(24 downto 0); 
    decim_35_q_fpga_out: out std_logic_vector(24 downto 0); 
    mix_i: out std_logic_vector(23 downto 0); 
    mix_q: out std_logic_vector(23 downto 0); 
    valid_f: out std_logic
  );
end channel2_tbt_entity_c5e2abdcfa;

architecture structural of channel2_tbt_entity_c5e2abdcfa is
  signal adc_ch2_i_net_x1: std_logic_vector(15 downto 0);
  signal ce_1_sg_x26: std_logic;
  signal ce_35_sg_x5: std_logic;
  signal ce_logic_1_sg_x14: std_logic;
  signal clk_1_sg_x26: std_logic;
  signal clk_35_sg_x5: std_logic;
  signal convert1_dout_net_x1: std_logic_vector(24 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(24 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x8: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x8: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x8: std_logic;
  signal delay6_q_net_x5: std_logic_vector(23 downto 0);
  signal delay7_q_net_x5: std_logic_vector(23 downto 0);
  signal fir_compiler_6_2_m_axis_data_tvalid_net_x0: std_logic;
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(24 downto 0);
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register5_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal register_q_net_x5: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);

begin
  adc_ch2_i_net_x1 <= adc_ch2_i;
  ce_1_sg_x26 <= ce_1;
  ce_35_sg_x5 <= ce_35;
  ce_logic_1_sg_x14 <= ce_logic_1;
  clk_1_sg_x26 <= clk_1;
  clk_35_sg_x5 <= clk_35;
  dds_m_axis_data_tdata_cosine_net_x8 <= dds_cosine_in;
  dds_m_axis_data_tdata_sine_net_x8 <= dds_msine_in;
  dds_m_axis_data_tvalid_net_x8 <= dds_valid_in;
  amp_f <= register5_q_net_x0;
  bpf_adc_fpga_out <= register_q_net_x5;
  decim_35_i_fpga_out <= convert2_dout_net_x1;
  decim_35_q_fpga_out <= convert1_dout_net_x1;
  mix_i <= delay7_q_net_x5;
  mix_q <= delay6_q_net_x5;
  valid_f <= register6_q_net_x0;

  ddc_1db418d5a4: entity work.ddc_entity_fbec30928b
    port map (
      adc_in => adc_ch2_i_net_x1,
      ce_1 => ce_1_sg_x26,
      ce_logic_1 => ce_logic_1_sg_x14,
      clk_1 => clk_1_sg_x26,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x8,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x8,
      dds_valid_in => dds_m_axis_data_tvalid_net_x8,
      bpf_out => register_q_net_x5,
      mix_i_out => delay7_q_net_x5,
      mix_q_out => delay6_q_net_x5
    );

  decim35_790814bb57: entity work.decim35_entity_3519cdb9ab
    port map (
      ce_1 => ce_1_sg_x26,
      ce_35 => ce_35_sg_x5,
      ce_logic_1 => ce_logic_1_sg_x14,
      clk_1 => clk_1_sg_x26,
      clk_35 => clk_35_sg_x5,
      i_in => delay7_q_net_x5,
      q_in => delay6_q_net_x5,
      i_out => convert2_dout_net_x1,
      q_out => convert1_dout_net_x1,
      valid_out => fir_compiler_6_2_m_axis_data_tvalid_net_x0
    );

  rect2pol: entity work.xlcordic_c062cc3a2d77ede2032de397150e15cd
    port map (
      ce => ce_35_sg_x5,
      clk => clk_35_sg_x5,
      s_axis_cartesian_tdata_imag => convert1_dout_net_x1,
      s_axis_cartesian_tdata_real => convert2_dout_net_x1,
      s_axis_cartesian_tvalid => fir_compiler_6_2_m_axis_data_tvalid_net_x0,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x5,
      clk => clk_35_sg_x5,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x5,
      clk => clk_35_sg_x5,
      d(0) => rect2pol_m_axis_dout_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Channel3_tbt"

entity channel3_tbt_entity_63129db436 is
  port (
    adc_ch3_i: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    ce_logic_1: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    dds_cosine_in: in std_logic_vector(23 downto 0); 
    dds_msine_in: in std_logic_vector(23 downto 0); 
    dds_valid_in: in std_logic; 
    amp_f: out std_logic_vector(24 downto 0); 
    bpf_adc_fpga_out: out std_logic_vector(23 downto 0); 
    decim_35_i_fpga_out: out std_logic_vector(24 downto 0); 
    decim_35_q_fpga_out: out std_logic_vector(24 downto 0); 
    mix_i: out std_logic_vector(23 downto 0); 
    mix_q: out std_logic_vector(23 downto 0); 
    valid_f: out std_logic
  );
end channel3_tbt_entity_63129db436;

architecture structural of channel3_tbt_entity_63129db436 is
  signal adc_ch3_i_net_x1: std_logic_vector(15 downto 0);
  signal ce_1_sg_x35: std_logic;
  signal ce_35_sg_x7: std_logic;
  signal ce_logic_1_sg_x19: std_logic;
  signal clk_1_sg_x35: std_logic;
  signal clk_35_sg_x7: std_logic;
  signal convert1_dout_net_x1: std_logic_vector(24 downto 0);
  signal convert2_dout_net_x1: std_logic_vector(24 downto 0);
  signal dds_m_axis_data_tdata_cosine_net_x11: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x11: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x11: std_logic;
  signal delay6_q_net_x5: std_logic_vector(23 downto 0);
  signal delay7_q_net_x5: std_logic_vector(23 downto 0);
  signal fir_compiler_6_2_m_axis_data_tvalid_net_x0: std_logic;
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(24 downto 0);
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register5_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal register_q_net_x5: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);

begin
  adc_ch3_i_net_x1 <= adc_ch3_i;
  ce_1_sg_x35 <= ce_1;
  ce_35_sg_x7 <= ce_35;
  ce_logic_1_sg_x19 <= ce_logic_1;
  clk_1_sg_x35 <= clk_1;
  clk_35_sg_x7 <= clk_35;
  dds_m_axis_data_tdata_cosine_net_x11 <= dds_cosine_in;
  dds_m_axis_data_tdata_sine_net_x11 <= dds_msine_in;
  dds_m_axis_data_tvalid_net_x11 <= dds_valid_in;
  amp_f <= register5_q_net_x0;
  bpf_adc_fpga_out <= register_q_net_x5;
  decim_35_i_fpga_out <= convert2_dout_net_x1;
  decim_35_q_fpga_out <= convert1_dout_net_x1;
  mix_i <= delay7_q_net_x5;
  mix_q <= delay6_q_net_x5;
  valid_f <= register6_q_net_x0;

  ddc_7682ff735a: entity work.ddc_entity_fbec30928b
    port map (
      adc_in => adc_ch3_i_net_x1,
      ce_1 => ce_1_sg_x35,
      ce_logic_1 => ce_logic_1_sg_x19,
      clk_1 => clk_1_sg_x35,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x11,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x11,
      dds_valid_in => dds_m_axis_data_tvalid_net_x11,
      bpf_out => register_q_net_x5,
      mix_i_out => delay7_q_net_x5,
      mix_q_out => delay6_q_net_x5
    );

  decim35_89edd3a010: entity work.decim35_entity_3519cdb9ab
    port map (
      ce_1 => ce_1_sg_x35,
      ce_35 => ce_35_sg_x7,
      ce_logic_1 => ce_logic_1_sg_x19,
      clk_1 => clk_1_sg_x35,
      clk_35 => clk_35_sg_x7,
      i_in => delay7_q_net_x5,
      q_in => delay6_q_net_x5,
      i_out => convert2_dout_net_x1,
      q_out => convert1_dout_net_x1,
      valid_out => fir_compiler_6_2_m_axis_data_tvalid_net_x0
    );

  rect2pol: entity work.xlcordic_c062cc3a2d77ede2032de397150e15cd
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      s_axis_cartesian_tdata_imag => convert1_dout_net_x1,
      s_axis_cartesian_tdata_real => convert2_dout_net_x1,
      s_axis_cartesian_tvalid => fir_compiler_6_2_m_axis_data_tvalid_net_x0,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d(0) => rect2pol_m_axis_dout_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Decim_Q_monit"

entity decim_q_monit_entity_d3ca57d66c is
  port (
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    ce_11130000: in std_logic; 
    ce_2782500: in std_logic; 
    ce_5565000: in std_logic; 
    ce_logic_1113: in std_logic; 
    ce_logic_2782500: in std_logic; 
    ce_logic_5565000: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    clk_11130000: in std_logic; 
    clk_2782500: in std_logic; 
    clk_5565000: in std_logic; 
    data_in: in std_logic_vector(23 downto 0); 
    monit_out: out std_logic_vector(23 downto 0)
  );
end decim_q_monit_entity_d3ca57d66c;

architecture structural of decim_q_monit_entity_d3ca57d66c is
  signal ce_11130000_sg_x0: std_logic;
  signal ce_1113_sg_x8: std_logic;
  signal ce_1_sg_x36: std_logic;
  signal ce_2782500_sg_x0: std_logic;
  signal ce_5565000_sg_x0: std_logic;
  signal ce_logic_1113_sg_x0: std_logic;
  signal ce_logic_2782500_sg_x0: std_logic;
  signal ce_logic_5565000_sg_x0: std_logic;
  signal cfir_monit_m_axis_data_tdata_net: std_logic_vector(40 downto 0);
  signal cfir_monit_m_axis_data_tvalid_net: std_logic;
  signal cic_monit_m_axis_data_tdata_data_net: std_logic_vector(23 downto 0);
  signal cic_monit_m_axis_data_tvalid_net: std_logic;
  signal clk_11130000_sg_x0: std_logic;
  signal clk_1113_sg_x8: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal clk_2782500_sg_x0: std_logic;
  signal clk_5565000_sg_x0: std_logic;
  signal convert1_dout_net: std_logic_vector(23 downto 0);
  signal convert2_dout_net: std_logic_vector(24 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal pfir_monit_m_axis_data_tdata_net: std_logic_vector(41 downto 0);
  signal pfir_monit_m_axis_data_tvalid_net: std_logic;
  signal register2_q_net: std_logic_vector(23 downto 0);
  signal register3_q_net: std_logic_vector(24 downto 0);
  signal register5_q_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x36 <= ce_1;
  ce_1113_sg_x8 <= ce_1113;
  ce_11130000_sg_x0 <= ce_11130000;
  ce_2782500_sg_x0 <= ce_2782500;
  ce_5565000_sg_x0 <= ce_5565000;
  ce_logic_1113_sg_x0 <= ce_logic_1113;
  ce_logic_2782500_sg_x0 <= ce_logic_2782500;
  ce_logic_5565000_sg_x0 <= ce_logic_5565000;
  clk_1_sg_x36 <= clk_1;
  clk_1113_sg_x8 <= clk_1113;
  clk_11130000_sg_x0 <= clk_11130000;
  clk_2782500_sg_x0 <= clk_2782500;
  clk_5565000_sg_x0 <= clk_5565000;
  down_sample2_q_net_x0 <= data_in;
  monit_out <= register5_q_net_x0;

  cfir_monit: entity work.xlfir_compiler_63d9ad3400f500cbd021770c26f451ad
    port map (
      ce => ce_1_sg_x36,
      ce_2782500 => ce_2782500_sg_x0,
      ce_5565000 => ce_5565000_sg_x0,
      ce_logic_2782500 => ce_logic_2782500_sg_x0,
      clk => clk_1_sg_x36,
      clk_2782500 => clk_2782500_sg_x0,
      clk_5565000 => clk_5565000_sg_x0,
      clk_logic_2782500 => clk_2782500_sg_x0,
      s_axis_data_tdata => register2_q_net,
      src_ce => ce_2782500_sg_x0,
      src_clk => clk_2782500_sg_x0,
      m_axis_data_tdata => cfir_monit_m_axis_data_tdata_net,
      m_axis_data_tvalid => cfir_monit_m_axis_data_tvalid_net
    );

  cic_monit: entity work.xlcic_compiler_95547d442151284e81277c01e1dd33ef
    port map (
      ce => ce_1_sg_x36,
      ce_1113 => ce_1113_sg_x8,
      ce_2782500 => ce_2782500_sg_x0,
      ce_logic_1113 => ce_logic_1113_sg_x0,
      clk => clk_1_sg_x36,
      clk_1113 => clk_1113_sg_x8,
      clk_2782500 => clk_2782500_sg_x0,
      clk_logic_1113 => clk_1113_sg_x8,
      s_axis_data_tdata_data => down_sample2_q_net_x0,
      m_axis_data_tdata_data => cic_monit_m_axis_data_tdata_data_net,
      m_axis_data_tvalid => cic_monit_m_axis_data_tvalid_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 38,
      din_width => 42,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_11130000_sg_x0,
      clk => clk_11130000_sg_x0,
      clr => '0',
      din => pfir_monit_m_axis_data_tdata_net,
      en => "1",
      dout => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 38,
      din_width => 41,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_5565000_sg_x0,
      clk => clk_5565000_sg_x0,
      clr => '0',
      din => cfir_monit_m_axis_data_tdata_net,
      en => "1",
      dout => convert2_dout_net
    );

  pfir_monit: entity work.xlfir_compiler_d0050991ffa08d9151315827675f900b
    port map (
      ce => ce_1_sg_x36,
      ce_11130000 => ce_11130000_sg_x0,
      ce_5565000 => ce_5565000_sg_x0,
      ce_logic_5565000 => ce_logic_5565000_sg_x0,
      clk => clk_1_sg_x36,
      clk_11130000 => clk_11130000_sg_x0,
      clk_5565000 => clk_5565000_sg_x0,
      clk_logic_5565000 => clk_5565000_sg_x0,
      s_axis_data_tdata => register3_q_net,
      src_ce => ce_5565000_sg_x0,
      src_clk => clk_5565000_sg_x0,
      m_axis_data_tdata => pfir_monit_m_axis_data_tdata_net,
      m_axis_data_tvalid => pfir_monit_m_axis_data_tvalid_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_2782500_sg_x0,
      clk => clk_2782500_sg_x0,
      d => reinterpret_output_port_net,
      en(0) => cic_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_5565000_sg_x0,
      clk => clk_5565000_sg_x0,
      d => convert2_dout_net,
      en(0) => cfir_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register3_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_11130000_sg_x0,
      clk => clk_11130000_sg_x0,
      d => convert1_dout_net,
      en(0) => pfir_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  reinterpret: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_monit_m_axis_data_tdata_data_net,
      output_port => reinterpret_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Decim_Sum_monit"

entity decim_sum_monit_entity_1ee5debdc8 is
  port (
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    ce_11130000: in std_logic; 
    ce_2782500: in std_logic; 
    ce_5565000: in std_logic; 
    ce_logic_1113: in std_logic; 
    ce_logic_2782500: in std_logic; 
    ce_logic_5565000: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    clk_11130000: in std_logic; 
    clk_2782500: in std_logic; 
    clk_5565000: in std_logic; 
    data_in: in std_logic_vector(23 downto 0); 
    monit_out: out std_logic_vector(23 downto 0)
  );
end decim_sum_monit_entity_1ee5debdc8;

architecture structural of decim_sum_monit_entity_1ee5debdc8 is
  signal ce_11130000_sg_x1: std_logic;
  signal ce_1113_sg_x9: std_logic;
  signal ce_1_sg_x37: std_logic;
  signal ce_2782500_sg_x1: std_logic;
  signal ce_5565000_sg_x1: std_logic;
  signal ce_logic_1113_sg_x1: std_logic;
  signal ce_logic_2782500_sg_x1: std_logic;
  signal ce_logic_5565000_sg_x1: std_logic;
  signal cfir_monit_m_axis_data_tdata_net: std_logic_vector(40 downto 0);
  signal cfir_monit_m_axis_data_tvalid_net: std_logic;
  signal cic_monit_m_axis_data_tdata_data_net: std_logic_vector(23 downto 0);
  signal cic_monit_m_axis_data_tvalid_net: std_logic;
  signal clk_11130000_sg_x1: std_logic;
  signal clk_1113_sg_x9: std_logic;
  signal clk_1_sg_x37: std_logic;
  signal clk_2782500_sg_x1: std_logic;
  signal clk_5565000_sg_x1: std_logic;
  signal convert1_dout_net: std_logic_vector(23 downto 0);
  signal convert2_dout_net: std_logic_vector(25 downto 0);
  signal down_sample3_q_net_x0: std_logic_vector(23 downto 0);
  signal pfir_monit_m_axis_data_tdata_net: std_logic_vector(42 downto 0);
  signal pfir_monit_m_axis_data_tvalid_net: std_logic;
  signal register2_q_net: std_logic_vector(23 downto 0);
  signal register3_q_net: std_logic_vector(25 downto 0);
  signal register5_q_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x37 <= ce_1;
  ce_1113_sg_x9 <= ce_1113;
  ce_11130000_sg_x1 <= ce_11130000;
  ce_2782500_sg_x1 <= ce_2782500;
  ce_5565000_sg_x1 <= ce_5565000;
  ce_logic_1113_sg_x1 <= ce_logic_1113;
  ce_logic_2782500_sg_x1 <= ce_logic_2782500;
  ce_logic_5565000_sg_x1 <= ce_logic_5565000;
  clk_1_sg_x37 <= clk_1;
  clk_1113_sg_x9 <= clk_1113;
  clk_11130000_sg_x1 <= clk_11130000;
  clk_2782500_sg_x1 <= clk_2782500;
  clk_5565000_sg_x1 <= clk_5565000;
  down_sample3_q_net_x0 <= data_in;
  monit_out <= register5_q_net_x0;

  cfir_monit: entity work.xlfir_compiler_8639b3660dc5b7c78f3b8f56b4679494
    port map (
      ce => ce_1_sg_x37,
      ce_2782500 => ce_2782500_sg_x1,
      ce_5565000 => ce_5565000_sg_x1,
      ce_logic_2782500 => ce_logic_2782500_sg_x1,
      clk => clk_1_sg_x37,
      clk_2782500 => clk_2782500_sg_x1,
      clk_5565000 => clk_5565000_sg_x1,
      clk_logic_2782500 => clk_2782500_sg_x1,
      s_axis_data_tdata => register2_q_net,
      src_ce => ce_2782500_sg_x1,
      src_clk => clk_2782500_sg_x1,
      m_axis_data_tdata => cfir_monit_m_axis_data_tdata_net,
      m_axis_data_tvalid => cfir_monit_m_axis_data_tvalid_net
    );

  cic_monit: entity work.xlcic_compiler_95547d442151284e81277c01e1dd33ef
    port map (
      ce => ce_1_sg_x37,
      ce_1113 => ce_1113_sg_x9,
      ce_2782500 => ce_2782500_sg_x1,
      ce_logic_1113 => ce_logic_1113_sg_x1,
      clk => clk_1_sg_x37,
      clk_1113 => clk_1113_sg_x9,
      clk_2782500 => clk_2782500_sg_x1,
      clk_logic_1113 => clk_1113_sg_x9,
      s_axis_data_tdata_data => down_sample3_q_net_x0,
      m_axis_data_tdata_data => cic_monit_m_axis_data_tdata_data_net,
      m_axis_data_tvalid => cic_monit_m_axis_data_tvalid_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 36,
      din_width => 43,
      dout_arith => 2,
      dout_bin_pt => 20,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_11130000_sg_x1,
      clk => clk_11130000_sg_x1,
      clr => '0',
      din => pfir_monit_m_axis_data_tdata_net,
      en => "1",
      dout => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 35,
      din_width => 41,
      dout_arith => 2,
      dout_bin_pt => 20,
      dout_width => 26,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_5565000_sg_x1,
      clk => clk_5565000_sg_x1,
      clr => '0',
      din => cfir_monit_m_axis_data_tdata_net,
      en => "1",
      dout => convert2_dout_net
    );

  pfir_monit: entity work.xlfir_compiler_472d6cb416f02569126e68c627373423
    port map (
      ce => ce_1_sg_x37,
      ce_11130000 => ce_11130000_sg_x1,
      ce_5565000 => ce_5565000_sg_x1,
      ce_logic_5565000 => ce_logic_5565000_sg_x1,
      clk => clk_1_sg_x37,
      clk_11130000 => clk_11130000_sg_x1,
      clk_5565000 => clk_5565000_sg_x1,
      clk_logic_5565000 => clk_5565000_sg_x1,
      s_axis_data_tdata => register3_q_net,
      src_ce => ce_5565000_sg_x1,
      src_clk => clk_5565000_sg_x1,
      m_axis_data_tdata => pfir_monit_m_axis_data_tdata_net,
      m_axis_data_tvalid => pfir_monit_m_axis_data_tvalid_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_2782500_sg_x1,
      clk => clk_2782500_sg_x1,
      d => reinterpret_output_port_net,
      en(0) => cic_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_5565000_sg_x1,
      clk => clk_5565000_sg_x1,
      d => convert2_dout_net,
      en(0) => cfir_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register3_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_11130000_sg_x1,
      clk => clk_11130000_sg_x1,
      d => convert1_dout_net,
      en(0) => pfir_monit_m_axis_data_tvalid_net,
      rst => "0",
      q => register5_q_net_x0
    );

  reinterpret: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_monit_m_axis_data_tdata_data_net,
      output_port => reinterpret_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb/DataReg_En"

entity datareg_en_entity_79473f9ed1 is
  port (
    ce_1113: in std_logic; 
    clk_1113: in std_logic; 
    din: in std_logic_vector(26 downto 0); 
    en: in std_logic; 
    dout: out std_logic_vector(26 downto 0)
  );
end datareg_en_entity_79473f9ed1;

architecture structural of datareg_en_entity_79473f9ed1 is
  signal ce_1113_sg_x12: std_logic;
  signal clk_1113_sg_x12: std_logic;
  signal delta_x_s_net_x0: std_logic_vector(26 downto 0);
  signal register17_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(26 downto 0);

begin
  ce_1113_sg_x12 <= ce_1113;
  clk_1113_sg_x12 <= clk_1113;
  delta_x_s_net_x0 <= din;
  register17_q_net_x0 <= en;
  dout <= register_q_net_x0;

  register_x0: entity work.xlregister
    generic map (
      d_width => 27,
      init_value => b"000000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x12,
      clk => clk_1113_sg_x12,
      d => delta_x_s_net_x0,
      en(0) => register17_q_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb/unsigned2signed1"

entity unsigned2signed1_entity_4871dec4a6 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    s_data: in std_logic_vector(26 downto 0); 
    u_data: in std_logic_vector(22 downto 0); 
    data_out: out std_logic_vector(23 downto 0)
  );
end unsigned2signed1_entity_4871dec4a6;

architecture structural of unsigned2signed1_entity_4871dec4a6 is
  signal ce_1_sg_x40: std_logic;
  signal clk_1_sg_x40: std_logic;
  signal concat_y_net: std_logic_vector(49 downto 0);
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(22 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(26 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(49 downto 0);
  signal y_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal y_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);

begin
  ce_1_sg_x40 <= ce_1;
  clk_1_sg_x40 <= clk_1;
  y_divider_m_axis_dout_tdata_quotient_net_x0 <= s_data;
  y_divider_m_axis_dout_tdata_fractional_net_x0 <= u_data;
  data_out <= convert_dout_net_x0;

  concat: entity work.concat_0d0fc5690d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret2_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 23,
      din_width => 50,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  reinterpret: entity work.reinterpret_1d284b35d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_48a79104f5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => y_divider_m_axis_dout_tdata_fractional_net_x0,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_bf9824e821
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => y_divider_m_axis_dout_tdata_quotient_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb"

entity delta_sigma_fofb_entity_ee61e649ea is
  port (
    a: in std_logic_vector(24 downto 0); 
    avalid: in std_logic; 
    b: in std_logic_vector(24 downto 0); 
    bvalid: in std_logic; 
    c: in std_logic_vector(24 downto 0); 
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    cvalid: in std_logic; 
    d: in std_logic_vector(24 downto 0); 
    delta_sigma_thres: in std_logic_vector(26 downto 0); 
    dvalid: in std_logic; 
    q: out std_logic_vector(23 downto 0); 
    sum_x0: out std_logic_vector(23 downto 0); 
    x: out std_logic_vector(23 downto 0); 
    y: out std_logic_vector(23 downto 0)
  );
end delta_sigma_fofb_entity_ee61e649ea;

architecture structural of delta_sigma_fofb_entity_ee61e649ea is
  signal a_plus_b_s_net: std_logic_vector(25 downto 0);
  signal a_plus_c_s_net: std_logic_vector(25 downto 0);
  signal a_plus_d_s_net: std_logic_vector(25 downto 0);
  signal b_plus_c_s_net: std_logic_vector(25 downto 0);
  signal b_plus_d_s_net: std_logic_vector(25 downto 0);
  signal c_plus_d_s_net: std_logic_vector(25 downto 0);
  signal ce_1113_sg_x16: std_logic;
  signal ce_1_sg_x43: std_logic;
  signal clk_1113_sg_x16: std_logic;
  signal clk_1_sg_x43: std_logic;
  signal convert_dout_net: std_logic_vector(23 downto 0);
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal convert_dout_net_x1: std_logic_vector(23 downto 0);
  signal convert_dout_net_x2: std_logic_vector(23 downto 0);
  signal del_sig_div_fofb_thres_i_net_x0: std_logic_vector(26 downto 0);
  signal delay_q_net: std_logic_vector(26 downto 0);
  signal delta_q_s_net_x0: std_logic_vector(26 downto 0);
  signal delta_x_s_net_x0: std_logic_vector(26 downto 0);
  signal delta_y_s_net_x0: std_logic_vector(26 downto 0);
  signal expression1_dout_net: std_logic;
  signal expression_dout_net: std_logic;
  signal fifo_q_dout_net: std_logic_vector(26 downto 0);
  signal fifo_q_empty_net: std_logic;
  signal fifo_sum_dout_net: std_logic_vector(26 downto 0);
  signal fifo_sum_empty_net: std_logic;
  signal fifo_x_dout_net: std_logic_vector(26 downto 0);
  signal fifo_x_empty_net: std_logic;
  signal fifo_y_dout_net: std_logic_vector(26 downto 0);
  signal fifo_y_empty_net: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal q_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal q_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal q_divider_m_axis_dout_tvalid_net: std_logic;
  signal q_divider_s_axis_dividend_tready_net: std_logic;
  signal q_divider_s_axis_divisor_tready_net: std_logic;
  signal register11_q_net_x0: std_logic_vector(23 downto 0);
  signal register12_q_net_x0: std_logic_vector(23 downto 0);
  signal register13_q_net_x0: std_logic_vector(23 downto 0);
  signal register17_q_net_x3: std_logic;
  signal register19_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(25 downto 0);
  signal register2_q_net: std_logic_vector(25 downto 0);
  signal register3_q_net: std_logic_vector(25 downto 0);
  signal register4_q_net: std_logic_vector(25 downto 0);
  signal register5_q_net: std_logic_vector(25 downto 0);
  signal register5_q_net_x4: std_logic_vector(24 downto 0);
  signal register5_q_net_x5: std_logic_vector(24 downto 0);
  signal register5_q_net_x6: std_logic_vector(24 downto 0);
  signal register5_q_net_x7: std_logic_vector(24 downto 0);
  signal register6_q_net: std_logic_vector(25 downto 0);
  signal register6_q_net_x4: std_logic;
  signal register6_q_net_x5: std_logic;
  signal register6_q_net_x6: std_logic;
  signal register6_q_net_x7: std_logic;
  signal register_q_net_x0: std_logic_vector(26 downto 0);
  signal register_q_net_x1: std_logic_vector(26 downto 0);
  signal register_q_net_x2: std_logic_vector(26 downto 0);
  signal register_q_net_x3: std_logic_vector(26 downto 0);
  signal relational_op_net: std_logic;
  signal sum_s_net_x0: std_logic_vector(26 downto 0);
  signal x_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal x_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal x_divider_m_axis_dout_tvalid_net: std_logic;
  signal x_divider_s_axis_dividend_tready_net: std_logic;
  signal x_divider_s_axis_divisor_tready_net: std_logic;
  signal y_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal y_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal y_divider_m_axis_dout_tvalid_net: std_logic;
  signal y_divider_s_axis_dividend_tready_net: std_logic;
  signal y_divider_s_axis_divisor_tready_net: std_logic;

begin
  register5_q_net_x4 <= a;
  register6_q_net_x4 <= avalid;
  register5_q_net_x5 <= b;
  register6_q_net_x5 <= bvalid;
  register5_q_net_x6 <= c;
  ce_1_sg_x43 <= ce_1;
  ce_1113_sg_x16 <= ce_1113;
  clk_1_sg_x43 <= clk_1;
  clk_1113_sg_x16 <= clk_1113;
  register6_q_net_x6 <= cvalid;
  register5_q_net_x7 <= d;
  del_sig_div_fofb_thres_i_net_x0 <= delta_sigma_thres;
  register6_q_net_x7 <= dvalid;
  q <= register12_q_net_x0;
  sum_x0 <= register19_q_net_x0;
  x <= register11_q_net_x0;
  y <= register13_q_net_x0;

  a_plus_b: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x5,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => a_plus_b_s_net
    );

  a_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x6,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => a_plus_c_s_net
    );

  a_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x7,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => a_plus_d_s_net
    );

  b_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x5,
      b => register5_q_net_x6,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => b_plus_c_s_net
    );

  b_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x5,
      b => register5_q_net_x7,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => b_plus_d_s_net
    );

  c_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x6,
      b => register5_q_net_x7,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => c_plus_d_s_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 23,
      din_width => 27,
      dout_arith => 2,
      dout_bin_pt => 20,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      din => delay_q_net,
      en => "1",
      dout => convert_dout_net
    );

  datareg_en1_3225c09afc: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1113 => ce_1113_sg_x16,
      clk_1113 => clk_1113_sg_x16,
      din => sum_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x1
    );

  datareg_en2_5b5f4b61b7: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1113 => ce_1113_sg_x16,
      clk_1113 => clk_1113_sg_x16,
      din => delta_y_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x2
    );

  datareg_en3_6643090018: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1113 => ce_1113_sg_x16,
      clk_1113 => clk_1113_sg_x16,
      din => delta_q_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x3
    );

  datareg_en_79473f9ed1: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1113 => ce_1113_sg_x16,
      clk_1113 => clk_1113_sg_x16,
      din => delta_x_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 39,
      reg_retiming => 0,
      reset => 0,
      width => 27
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => fifo_sum_dout_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delta_q: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register5_q_net,
      b => register6_q_net,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => delta_q_s_net_x0
    );

  delta_x: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register1_q_net,
      b => register3_q_net,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => delta_x_s_net_x0
    );

  delta_y: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register2_q_net,
      b => register4_q_net,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => delta_y_s_net_x0
    );

  expression: entity work.expr_24cbf78c62
    port map (
      a(0) => register6_q_net_x4,
      b(0) => register6_q_net_x5,
      c(0) => register6_q_net_x6,
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => register6_q_net_x7,
      dout(0) => expression_dout_net
    );

  expression1: entity work.expr_375d7bbece
    port map (
      a(0) => x_divider_s_axis_divisor_tready_net,
      b(0) => y_divider_s_axis_divisor_tready_net,
      c(0) => q_divider_s_axis_divisor_tready_net,
      ce => '0',
      clk => '0',
      clr => '0',
      dout(0) => expression1_dout_net
    );

  fifo_q: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      din => register_q_net_x3,
      en => '1',
      re => q_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x43,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x43,
      dout => fifo_q_dout_net,
      empty => fifo_q_empty_net
    );

  fifo_sum: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      din => register_q_net_x1,
      en => '1',
      re => expression1_dout_net,
      re_ce => ce_1_sg_x43,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x43,
      dout => fifo_sum_dout_net,
      empty => fifo_sum_empty_net
    );

  fifo_x: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      din => register_q_net_x0,
      en => '1',
      re => x_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x43,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x43,
      dout => fifo_x_dout_net,
      empty => fifo_x_empty_net
    );

  fifo_y: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      din => register_q_net_x2,
      en => '1',
      re => y_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x43,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x43,
      dout => fifo_y_dout_net,
      empty => fifo_y_empty_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip(0) => fifo_x_empty_net,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip(0) => fifo_sum_empty_net,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip(0) => fifo_y_empty_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip(0) => fifo_q_empty_net,
      op(0) => inverter3_op_net
    );

  q_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      s_axis_dividend_tdata_dividend => fifo_q_dout_net,
      s_axis_dividend_tvalid => inverter3_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => q_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => q_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => q_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => q_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => q_divider_s_axis_divisor_tready_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => b_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register11: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => convert_dout_net_x1,
      en(0) => x_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register11_q_net_x0
    );

  register12: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => convert_dout_net_x2,
      en(0) => q_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register12_q_net_x0
    );

  register13: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => convert_dout_net_x0,
      en(0) => y_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register13_q_net_x0
    );

  register17: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d(0) => expression_dout_net,
      en => "1",
      rst => "0",
      q(0) => register17_q_net_x3
    );

  register19: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d => convert_dout_net,
      en => "1",
      rst => "0",
      q => register19_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => a_plus_b_s_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => a_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => c_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => a_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      d => b_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register6_q_net
    );

  relational: entity work.relational_6505656e93
    port map (
      a => register_q_net_x1,
      b => del_sig_div_fofb_thres_i_net_x0,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  sum: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_2f1626aeedb3c308",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register3_q_net,
      b => register1_q_net,
      ce => ce_1113_sg_x16,
      clk => clk_1113_sg_x16,
      clr => '0',
      en => "1",
      s => sum_s_net_x0
    );

  unsigned2signed1_4871dec4a6: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x43,
      clk_1 => clk_1_sg_x43,
      s_data => y_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => y_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x0
    );

  unsigned2signed2_2f05b465d2: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x43,
      clk_1 => clk_1_sg_x43,
      s_data => x_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => x_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x1
    );

  unsigned2signed3_5318c8a639: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x43,
      clk_1 => clk_1_sg_x43,
      s_data => q_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => q_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x2
    );

  x_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      s_axis_dividend_tdata_dividend => fifo_x_dout_net,
      s_axis_dividend_tvalid => inverter_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => x_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => x_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => x_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => x_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => x_divider_s_axis_divisor_tready_net
    );

  y_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      s_axis_dividend_tdata_dividend => fifo_y_dout_net,
      s_axis_dividend_tvalid => inverter2_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => y_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => y_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => y_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => y_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => y_divider_s_axis_divisor_tready_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_tbt/DataReg_En"

entity datareg_en_entity_ed948c360a is
  port (
    ce_35: in std_logic; 
    clk_35: in std_logic; 
    din: in std_logic_vector(26 downto 0); 
    en: in std_logic; 
    dout: out std_logic_vector(26 downto 0)
  );
end datareg_en_entity_ed948c360a;

architecture structural of datareg_en_entity_ed948c360a is
  signal ce_35_sg_x8: std_logic;
  signal clk_35_sg_x8: std_logic;
  signal delta_x_s_net_x0: std_logic_vector(26 downto 0);
  signal register17_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(26 downto 0);

begin
  ce_35_sg_x8 <= ce_35;
  clk_35_sg_x8 <= clk_35;
  delta_x_s_net_x0 <= din;
  register17_q_net_x0 <= en;
  dout <= register_q_net_x0;

  register_x0: entity work.xlregister
    generic map (
      d_width => 27,
      init_value => b"000000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x8,
      clk => clk_35_sg_x8,
      d => delta_x_s_net_x0,
      en(0) => register17_q_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_tbt"

entity delta_sigma_tbt_entity_bbfa8a8a69 is
  port (
    a: in std_logic_vector(24 downto 0); 
    avalid: in std_logic; 
    b: in std_logic_vector(24 downto 0); 
    bvalid: in std_logic; 
    c: in std_logic_vector(24 downto 0); 
    ce_1: in std_logic; 
    ce_35: in std_logic; 
    clk_1: in std_logic; 
    clk_35: in std_logic; 
    cvalid: in std_logic; 
    d: in std_logic_vector(24 downto 0); 
    delta_sigma_thres: in std_logic_vector(26 downto 0); 
    dvalid: in std_logic; 
    q: out std_logic_vector(23 downto 0); 
    sum_x0: out std_logic_vector(23 downto 0); 
    x: out std_logic_vector(23 downto 0); 
    y: out std_logic_vector(23 downto 0)
  );
end delta_sigma_tbt_entity_bbfa8a8a69;

architecture structural of delta_sigma_tbt_entity_bbfa8a8a69 is
  signal a_plus_b_s_net: std_logic_vector(25 downto 0);
  signal a_plus_c_s_net: std_logic_vector(25 downto 0);
  signal a_plus_d_s_net: std_logic_vector(25 downto 0);
  signal b_plus_c_s_net: std_logic_vector(25 downto 0);
  signal b_plus_d_s_net: std_logic_vector(25 downto 0);
  signal c_plus_d_s_net: std_logic_vector(25 downto 0);
  signal ce_1_sg_x47: std_logic;
  signal ce_35_sg_x12: std_logic;
  signal clk_1_sg_x47: std_logic;
  signal clk_35_sg_x12: std_logic;
  signal convert_dout_net: std_logic_vector(23 downto 0);
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal convert_dout_net_x1: std_logic_vector(23 downto 0);
  signal convert_dout_net_x2: std_logic_vector(23 downto 0);
  signal del_sig_div_tbt_thres_i_net_x0: std_logic_vector(26 downto 0);
  signal delay_q_net: std_logic_vector(26 downto 0);
  signal delta_q_s_net_x0: std_logic_vector(26 downto 0);
  signal delta_x_s_net_x0: std_logic_vector(26 downto 0);
  signal delta_y_s_net_x0: std_logic_vector(26 downto 0);
  signal expression1_dout_net: std_logic;
  signal expression_dout_net: std_logic;
  signal fifo_q_dout_net: std_logic_vector(26 downto 0);
  signal fifo_q_empty_net: std_logic;
  signal fifo_sum_dout_net: std_logic_vector(26 downto 0);
  signal fifo_sum_empty_net: std_logic;
  signal fifo_x_dout_net: std_logic_vector(26 downto 0);
  signal fifo_x_empty_net: std_logic;
  signal fifo_y_dout_net: std_logic_vector(26 downto 0);
  signal fifo_y_empty_net: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal q_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal q_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal q_divider_m_axis_dout_tvalid_net: std_logic;
  signal q_divider_s_axis_dividend_tready_net: std_logic;
  signal q_divider_s_axis_divisor_tready_net: std_logic;
  signal register11_q_net_x0: std_logic_vector(23 downto 0);
  signal register12_q_net_x0: std_logic_vector(23 downto 0);
  signal register13_q_net_x0: std_logic_vector(23 downto 0);
  signal register17_q_net_x3: std_logic;
  signal register19_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(25 downto 0);
  signal register2_q_net: std_logic_vector(25 downto 0);
  signal register3_q_net: std_logic_vector(25 downto 0);
  signal register4_q_net: std_logic_vector(25 downto 0);
  signal register5_q_net: std_logic_vector(25 downto 0);
  signal register5_q_net_x4: std_logic_vector(24 downto 0);
  signal register5_q_net_x5: std_logic_vector(24 downto 0);
  signal register5_q_net_x6: std_logic_vector(24 downto 0);
  signal register5_q_net_x7: std_logic_vector(24 downto 0);
  signal register6_q_net: std_logic_vector(25 downto 0);
  signal register6_q_net_x4: std_logic;
  signal register6_q_net_x5: std_logic;
  signal register6_q_net_x6: std_logic;
  signal register6_q_net_x7: std_logic;
  signal register_q_net_x0: std_logic_vector(26 downto 0);
  signal register_q_net_x1: std_logic_vector(26 downto 0);
  signal register_q_net_x2: std_logic_vector(26 downto 0);
  signal register_q_net_x3: std_logic_vector(26 downto 0);
  signal relational_op_net: std_logic;
  signal sum_s_net_x0: std_logic_vector(26 downto 0);
  signal x_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal x_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal x_divider_m_axis_dout_tvalid_net: std_logic;
  signal x_divider_s_axis_dividend_tready_net: std_logic;
  signal x_divider_s_axis_divisor_tready_net: std_logic;
  signal y_divider_m_axis_dout_tdata_fractional_net_x0: std_logic_vector(22 downto 0);
  signal y_divider_m_axis_dout_tdata_quotient_net_x0: std_logic_vector(26 downto 0);
  signal y_divider_m_axis_dout_tvalid_net: std_logic;
  signal y_divider_s_axis_dividend_tready_net: std_logic;
  signal y_divider_s_axis_divisor_tready_net: std_logic;

begin
  register5_q_net_x4 <= a;
  register6_q_net_x4 <= avalid;
  register5_q_net_x5 <= b;
  register6_q_net_x5 <= bvalid;
  register5_q_net_x6 <= c;
  ce_1_sg_x47 <= ce_1;
  ce_35_sg_x12 <= ce_35;
  clk_1_sg_x47 <= clk_1;
  clk_35_sg_x12 <= clk_35;
  register6_q_net_x6 <= cvalid;
  register5_q_net_x7 <= d;
  del_sig_div_tbt_thres_i_net_x0 <= delta_sigma_thres;
  register6_q_net_x7 <= dvalid;
  q <= register12_q_net_x0;
  sum_x0 <= register19_q_net_x0;
  x <= register11_q_net_x0;
  y <= register13_q_net_x0;

  a_plus_b: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x5,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => a_plus_b_s_net
    );

  a_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x6,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => a_plus_c_s_net
    );

  a_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x4,
      b => register5_q_net_x7,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => a_plus_d_s_net
    );

  b_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x5,
      b => register5_q_net_x6,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => b_plus_c_s_net
    );

  b_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x5,
      b => register5_q_net_x7,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => b_plus_d_s_net
    );

  c_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_239e4f614ba09ab1",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 26
    )
    port map (
      a => register5_q_net_x6,
      b => register5_q_net_x7,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => c_plus_d_s_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 23,
      din_width => 27,
      dout_arith => 2,
      dout_bin_pt => 20,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      din => delay_q_net,
      en => "1",
      dout => convert_dout_net
    );

  datareg_en1_e5d0399944: entity work.datareg_en_entity_ed948c360a
    port map (
      ce_35 => ce_35_sg_x12,
      clk_35 => clk_35_sg_x12,
      din => sum_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x1
    );

  datareg_en2_02a2053e69: entity work.datareg_en_entity_ed948c360a
    port map (
      ce_35 => ce_35_sg_x12,
      clk_35 => clk_35_sg_x12,
      din => delta_y_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x2
    );

  datareg_en3_78179f99cc: entity work.datareg_en_entity_ed948c360a
    port map (
      ce_35 => ce_35_sg_x12,
      clk_35 => clk_35_sg_x12,
      din => delta_q_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x3
    );

  datareg_en_ed948c360a: entity work.datareg_en_entity_ed948c360a
    port map (
      ce_35 => ce_35_sg_x12,
      clk_35 => clk_35_sg_x12,
      din => delta_x_s_net_x0,
      en => register17_q_net_x3,
      dout => register_q_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 29,
      reg_retiming => 0,
      reset => 0,
      width => 27
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => fifo_sum_dout_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delta_q: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register5_q_net,
      b => register6_q_net,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => delta_q_s_net_x0
    );

  delta_x: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register1_q_net,
      b => register3_q_net,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => delta_x_s_net_x0
    );

  delta_y: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_1482f9e8df81448a",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register2_q_net,
      b => register4_q_net,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => delta_y_s_net_x0
    );

  expression: entity work.expr_24cbf78c62
    port map (
      a(0) => register6_q_net_x4,
      b(0) => register6_q_net_x5,
      c(0) => register6_q_net_x6,
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => register6_q_net_x7,
      dout(0) => expression_dout_net
    );

  expression1: entity work.expr_375d7bbece
    port map (
      a(0) => x_divider_s_axis_divisor_tready_net,
      b(0) => y_divider_s_axis_divisor_tready_net,
      c(0) => q_divider_s_axis_divisor_tready_net,
      ce => '0',
      clk => '0',
      clr => '0',
      dout(0) => expression1_dout_net
    );

  fifo_q: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      din => register_q_net_x3,
      en => '1',
      re => q_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x47,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x47,
      dout => fifo_q_dout_net,
      empty => fifo_q_empty_net
    );

  fifo_sum: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      din => register_q_net_x1,
      en => '1',
      re => expression1_dout_net,
      re_ce => ce_1_sg_x47,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x47,
      dout => fifo_sum_dout_net,
      empty => fifo_sum_empty_net
    );

  fifo_x: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      din => register_q_net_x0,
      en => '1',
      re => x_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x47,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x47,
      dout => fifo_x_dout_net,
      empty => fifo_x_empty_net
    );

  fifo_y: entity work.xlfifogen
    generic map (
      core_name0 => "fifo_fg84_26bc5f646d342e7f",
      data_count_width => 7,
      data_width => 27,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      din => register_q_net_x2,
      en => '1',
      re => y_divider_s_axis_dividend_tready_net,
      re_ce => ce_1_sg_x47,
      rst => '1',
      we => relational_op_net,
      we_ce => ce_1_sg_x47,
      dout => fifo_y_dout_net,
      empty => fifo_y_empty_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      ip(0) => fifo_x_empty_net,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      ip(0) => fifo_sum_empty_net,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      ip(0) => fifo_y_empty_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      clr => '0',
      ip(0) => fifo_q_empty_net,
      op(0) => inverter3_op_net
    );

  q_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      s_axis_dividend_tdata_dividend => fifo_q_dout_net,
      s_axis_dividend_tvalid => inverter3_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => q_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => q_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => q_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => q_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => q_divider_s_axis_divisor_tready_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => b_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register11: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => convert_dout_net_x1,
      en(0) => x_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register11_q_net_x0
    );

  register12: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => convert_dout_net_x2,
      en(0) => q_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register12_q_net_x0
    );

  register13: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => convert_dout_net_x0,
      en(0) => y_divider_m_axis_dout_tvalid_net,
      rst => "0",
      q => register13_q_net_x0
    );

  register17: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d(0) => expression_dout_net,
      en => "1",
      rst => "0",
      q(0) => register17_q_net_x3
    );

  register19: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => convert_dout_net,
      en => "1",
      rst => "0",
      q => register19_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => a_plus_b_s_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => a_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => c_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => a_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => b_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register6_q_net
    );

  relational: entity work.relational_6505656e93
    port map (
      a => register_q_net_x1,
      b => del_sig_div_tbt_thres_i_net_x0,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  sum: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 23,
      a_width => 26,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 26,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 27,
      core_name0 => "addsb_11_0_2f1626aeedb3c308",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 27,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 23,
      s_width => 27
    )
    port map (
      a => register3_q_net,
      b => register1_q_net,
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      clr => '0',
      en => "1",
      s => sum_s_net_x0
    );

  unsigned2signed1_0c64554e20: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x47,
      clk_1 => clk_1_sg_x47,
      s_data => y_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => y_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x0
    );

  unsigned2signed2_b5112b4796: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x47,
      clk_1 => clk_1_sg_x47,
      s_data => x_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => x_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x1
    );

  unsigned2signed3_3e8ecc04fc: entity work.unsigned2signed1_entity_4871dec4a6
    port map (
      ce_1 => ce_1_sg_x47,
      clk_1 => clk_1_sg_x47,
      s_data => q_divider_m_axis_dout_tdata_quotient_net_x0,
      u_data => q_divider_m_axis_dout_tdata_fractional_net_x0,
      data_out => convert_dout_net_x2
    );

  x_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      s_axis_dividend_tdata_dividend => fifo_x_dout_net,
      s_axis_dividend_tvalid => inverter_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => x_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => x_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => x_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => x_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => x_divider_s_axis_divisor_tready_net
    );

  y_divider: entity work.xldivider_generator_abfd96133d2f7eb1baefa6637fb34af7
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      s_axis_dividend_tdata_dividend => fifo_y_dout_net,
      s_axis_dividend_tvalid => inverter2_op_net,
      s_axis_divisor_tdata_divisor => fifo_sum_dout_net,
      s_axis_divisor_tvalid => inverter1_op_net,
      m_axis_dout_tdata_fractional => y_divider_m_axis_dout_tdata_fractional_net_x0,
      m_axis_dout_tdata_quotient => y_divider_m_axis_dout_tdata_quotient_net_x0,
      m_axis_dout_tvalid => y_divider_m_axis_dout_tvalid_net,
      s_axis_dividend_tready => y_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => y_divider_s_axis_divisor_tready_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066"

entity ddc_bpm_476_066 is
  port (
    adc_ch0_i: in std_logic_vector(15 downto 0); 
    adc_ch1_i: in std_logic_vector(15 downto 0); 
    adc_ch2_i: in std_logic_vector(15 downto 0); 
    adc_ch3_i: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    ce_1113: in std_logic; 
    ce_11130000: in std_logic; 
    ce_2782500: in std_logic; 
    ce_35: in std_logic; 
    ce_5565000: in std_logic; 
    ce_logic_1: in std_logic; 
    ce_logic_1113: in std_logic; 
    ce_logic_2782500: in std_logic; 
    ce_logic_5565000: in std_logic; 
    clk_1: in std_logic; 
    clk_1113: in std_logic; 
    clk_11130000: in std_logic; 
    clk_2782500: in std_logic; 
    clk_35: in std_logic; 
    clk_5565000: in std_logic; 
    del_sig_div_fofb_thres_i: in std_logic_vector(26 downto 0); 
    del_sig_div_tbt_thres_i: in std_logic_vector(26 downto 0); 
    adc_ch0_dbg_data_o: out std_logic_vector(15 downto 0); 
    adc_ch1_dbg_data_o: out std_logic_vector(15 downto 0); 
    adc_ch2_dbg_data_o: out std_logic_vector(15 downto 0); 
    adc_ch3_dbg_data_o: out std_logic_vector(15 downto 0); 
    bpf_ch0_o: out std_logic_vector(23 downto 0); 
    bpf_ch1_o: out std_logic_vector(23 downto 0); 
    bpf_ch2_o: out std_logic_vector(23 downto 0); 
    bpf_ch3_o: out std_logic_vector(23 downto 0); 
    cic_fofb_ch0_i_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch0_q_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch1_i_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch1_q_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch2_i_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch2_q_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch3_i_o: out std_logic_vector(24 downto 0); 
    cic_fofb_ch3_q_o: out std_logic_vector(24 downto 0); 
    fofb_amp_ch0_o: out std_logic_vector(24 downto 0); 
    fofb_amp_ch1_o: out std_logic_vector(24 downto 0); 
    fofb_amp_ch2_o: out std_logic_vector(24 downto 0); 
    fofb_amp_ch3_o: out std_logic_vector(24 downto 0); 
    mix_ch0_i_o: out std_logic_vector(23 downto 0); 
    mix_ch0_q_o: out std_logic_vector(23 downto 0); 
    mix_ch1_i_o: out std_logic_vector(23 downto 0); 
    mix_ch1_q_o: out std_logic_vector(23 downto 0); 
    mix_ch2_i_o: out std_logic_vector(23 downto 0); 
    mix_ch2_q_o: out std_logic_vector(23 downto 0); 
    mix_ch3_i_o: out std_logic_vector(23 downto 0); 
    mix_ch3_q_o: out std_logic_vector(23 downto 0); 
    poly35_ch0_i_o: out std_logic_vector(24 downto 0); 
    poly35_ch0_q_o: out std_logic_vector(24 downto 0); 
    poly35_ch1_i_o: out std_logic_vector(24 downto 0); 
    poly35_ch1_q_o: out std_logic_vector(24 downto 0); 
    poly35_ch2_i_o: out std_logic_vector(24 downto 0); 
    poly35_ch2_q_o: out std_logic_vector(24 downto 0); 
    poly35_ch3_i_o: out std_logic_vector(24 downto 0); 
    poly35_ch3_q_o: out std_logic_vector(24 downto 0); 
    q_fofb_o: out std_logic_vector(23 downto 0); 
    q_monit_o: out std_logic_vector(23 downto 0); 
    q_tbt_o: out std_logic_vector(23 downto 0); 
    sum_fofb_o: out std_logic_vector(23 downto 0); 
    sum_monit_o: out std_logic_vector(23 downto 0); 
    sum_tbt_o: out std_logic_vector(23 downto 0); 
    tbt_amp_ch0_o: out std_logic_vector(24 downto 0); 
    tbt_amp_ch1_o: out std_logic_vector(24 downto 0); 
    tbt_amp_ch2_o: out std_logic_vector(24 downto 0); 
    tbt_amp_ch3_o: out std_logic_vector(24 downto 0); 
    x_fofb_o: out std_logic_vector(23 downto 0); 
    x_monit_o: out std_logic_vector(23 downto 0); 
    x_tbt_o: out std_logic_vector(23 downto 0); 
    y_fofb_o: out std_logic_vector(23 downto 0); 
    y_monit_o: out std_logic_vector(23 downto 0); 
    y_tbt_o: out std_logic_vector(23 downto 0)
  );
end ddc_bpm_476_066;

architecture structural of ddc_bpm_476_066 is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "ddc_bpm_476_066,sysgen_core,{clock_period=8.88232184,clocking=Clock_Enables,compilation=HDL_Netlist,sample_periods=1.00000000000 35.00000000000 1113.00000000000 2782500.00000000000 5565000.00000000000 11130000.00000000000,testbench=0,total_blocks=1452,xilinx_adder_subtracter_block=20,xilinx_arithmetic_relational_operator_block=2,xilinx_bitwise_expression_evaluator_block=4,xilinx_bus_concatenator_block=6,xilinx_cic_compiler_3_0_block=12,xilinx_clock_enable_probe_block=3,xilinx_complex_multiplier_5_0__block=4,xilinx_constant_block_block=9,xilinx_cordic_5_0_block=8,xilinx_dds_compiler_5_0_block=1,xilinx_delay_block=26,xilinx_divider_generator_4_0_block=6,xilinx_down_sampler_block=4,xilinx_fifo_block_block=8,xilinx_fir_compiler_6_2_block=4,xilinx_fir_compiler_6_3_block=12,xilinx_gateway_in_block=6,xilinx_gateway_out_block=155,xilinx_inverter_block=8,xilinx_register_block=106,xilinx_sample_time_block_block=12,xilinx_system_generator_block=1,xilinx_type_converter_block=36,xilinx_type_reinterpreter_block=62,}";

  signal adc_ch0_i_net_x2: std_logic_vector(15 downto 0);
  signal adc_ch1_i_net_x2: std_logic_vector(15 downto 0);
  signal adc_ch2_i_net_x2: std_logic_vector(15 downto 0);
  signal adc_ch3_i_net_x2: std_logic_vector(15 downto 0);
  signal bpf_ch0_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch1_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch2_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch3_o_net: std_logic_vector(23 downto 0);
  signal ce_11130000_sg_x4: std_logic;
  signal ce_1113_sg_x17: std_logic;
  signal ce_1_sg_x48: std_logic;
  signal ce_2782500_sg_x4: std_logic;
  signal ce_35_sg_x13: std_logic;
  signal ce_5565000_sg_x4: std_logic;
  signal ce_logic_1113_sg_x4: std_logic;
  signal ce_logic_1_sg_x20: std_logic;
  signal ce_logic_2782500_sg_x4: std_logic;
  signal ce_logic_5565000_sg_x4: std_logic;
  signal cic_fofb_ch0_i_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch0_q_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch1_i_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch1_q_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch2_i_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch2_q_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch3_i_o_net: std_logic_vector(24 downto 0);
  signal cic_fofb_ch3_q_o_net: std_logic_vector(24 downto 0);
  signal clk_11130000_sg_x4: std_logic;
  signal clk_1113_sg_x17: std_logic;
  signal clk_1_sg_x48: std_logic;
  signal clk_2782500_sg_x4: std_logic;
  signal clk_35_sg_x13: std_logic;
  signal clk_5565000_sg_x4: std_logic;
  signal constant3_op_net: std_logic;
  signal dds_m_axis_data_tdata_cosine_net_x11: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tdata_sine_net_x11: std_logic_vector(23 downto 0);
  signal dds_m_axis_data_tvalid_net_x11: std_logic;
  signal del_sig_div_fofb_thres_i_net: std_logic_vector(26 downto 0);
  signal del_sig_div_tbt_thres_i_net: std_logic_vector(26 downto 0);
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(23 downto 0);
  signal fofb_amp_ch0_o_net: std_logic_vector(24 downto 0);
  signal fofb_amp_ch1_o_net: std_logic_vector(24 downto 0);
  signal fofb_amp_ch2_o_net: std_logic_vector(24 downto 0);
  signal fofb_amp_ch3_o_net: std_logic_vector(24 downto 0);
  signal mix_ch0_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch0_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch1_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch1_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch2_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch2_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch3_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch3_q_o_net: std_logic_vector(23 downto 0);
  signal poly35_ch0_i_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch0_q_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch1_i_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch1_q_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch2_i_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch2_q_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch3_i_o_net: std_logic_vector(24 downto 0);
  signal poly35_ch3_q_o_net: std_logic_vector(24 downto 0);
  signal q_fofb_o_net: std_logic_vector(23 downto 0);
  signal q_monit_o_net: std_logic_vector(23 downto 0);
  signal q_tbt_o_net: std_logic_vector(23 downto 0);
  signal register6_q_net_x10: std_logic;
  signal register6_q_net_x11: std_logic;
  signal register6_q_net_x4: std_logic;
  signal register6_q_net_x5: std_logic;
  signal register6_q_net_x6: std_logic;
  signal register6_q_net_x7: std_logic;
  signal register6_q_net_x8: std_logic;
  signal register6_q_net_x9: std_logic;
  signal sum_fofb_o_net: std_logic_vector(23 downto 0);
  signal sum_monit_o_net: std_logic_vector(23 downto 0);
  signal sum_tbt_o_net: std_logic_vector(23 downto 0);
  signal tbt_amp_ch0_o_net: std_logic_vector(24 downto 0);
  signal tbt_amp_ch1_o_net: std_logic_vector(24 downto 0);
  signal tbt_amp_ch2_o_net: std_logic_vector(24 downto 0);
  signal tbt_amp_ch3_o_net: std_logic_vector(24 downto 0);
  signal x_fofb_o_net: std_logic_vector(23 downto 0);
  signal x_monit_o_net: std_logic_vector(23 downto 0);
  signal x_tbt_o_net: std_logic_vector(23 downto 0);
  signal y_fofb_o_net: std_logic_vector(23 downto 0);
  signal y_monit_o_net: std_logic_vector(23 downto 0);
  signal y_tbt_o_net: std_logic_vector(23 downto 0);

begin
  adc_ch0_i_net_x2 <= adc_ch0_i;
  adc_ch1_i_net_x2 <= adc_ch1_i;
  adc_ch2_i_net_x2 <= adc_ch2_i;
  adc_ch3_i_net_x2 <= adc_ch3_i;
  ce_1_sg_x48 <= ce_1;
  ce_1113_sg_x17 <= ce_1113;
  ce_11130000_sg_x4 <= ce_11130000;
  ce_2782500_sg_x4 <= ce_2782500;
  ce_35_sg_x13 <= ce_35;
  ce_5565000_sg_x4 <= ce_5565000;
  ce_logic_1_sg_x20 <= ce_logic_1;
  ce_logic_1113_sg_x4 <= ce_logic_1113;
  ce_logic_2782500_sg_x4 <= ce_logic_2782500;
  ce_logic_5565000_sg_x4 <= ce_logic_5565000;
  clk_1_sg_x48 <= clk_1;
  clk_1113_sg_x17 <= clk_1113;
  clk_11130000_sg_x4 <= clk_11130000;
  clk_2782500_sg_x4 <= clk_2782500;
  clk_35_sg_x13 <= clk_35;
  clk_5565000_sg_x4 <= clk_5565000;
  del_sig_div_fofb_thres_i_net <= del_sig_div_fofb_thres_i;
  del_sig_div_tbt_thres_i_net <= del_sig_div_tbt_thres_i;
  adc_ch0_dbg_data_o <= adc_ch0_i_net_x2;
  adc_ch1_dbg_data_o <= adc_ch1_i_net_x2;
  adc_ch2_dbg_data_o <= adc_ch2_i_net_x2;
  adc_ch3_dbg_data_o <= adc_ch3_i_net_x2;
  bpf_ch0_o <= bpf_ch0_o_net;
  bpf_ch1_o <= bpf_ch1_o_net;
  bpf_ch2_o <= bpf_ch2_o_net;
  bpf_ch3_o <= bpf_ch3_o_net;
  cic_fofb_ch0_i_o <= cic_fofb_ch0_i_o_net;
  cic_fofb_ch0_q_o <= cic_fofb_ch0_q_o_net;
  cic_fofb_ch1_i_o <= cic_fofb_ch1_i_o_net;
  cic_fofb_ch1_q_o <= cic_fofb_ch1_q_o_net;
  cic_fofb_ch2_i_o <= cic_fofb_ch2_i_o_net;
  cic_fofb_ch2_q_o <= cic_fofb_ch2_q_o_net;
  cic_fofb_ch3_i_o <= cic_fofb_ch3_i_o_net;
  cic_fofb_ch3_q_o <= cic_fofb_ch3_q_o_net;
  fofb_amp_ch0_o <= fofb_amp_ch0_o_net;
  fofb_amp_ch1_o <= fofb_amp_ch1_o_net;
  fofb_amp_ch2_o <= fofb_amp_ch2_o_net;
  fofb_amp_ch3_o <= fofb_amp_ch3_o_net;
  mix_ch0_i_o <= mix_ch0_i_o_net;
  mix_ch0_q_o <= mix_ch0_q_o_net;
  mix_ch1_i_o <= mix_ch1_i_o_net;
  mix_ch1_q_o <= mix_ch1_q_o_net;
  mix_ch2_i_o <= mix_ch2_i_o_net;
  mix_ch2_q_o <= mix_ch2_q_o_net;
  mix_ch3_i_o <= mix_ch3_i_o_net;
  mix_ch3_q_o <= mix_ch3_q_o_net;
  poly35_ch0_i_o <= poly35_ch0_i_o_net;
  poly35_ch0_q_o <= poly35_ch0_q_o_net;
  poly35_ch1_i_o <= poly35_ch1_i_o_net;
  poly35_ch1_q_o <= poly35_ch1_q_o_net;
  poly35_ch2_i_o <= poly35_ch2_i_o_net;
  poly35_ch2_q_o <= poly35_ch2_q_o_net;
  poly35_ch3_i_o <= poly35_ch3_i_o_net;
  poly35_ch3_q_o <= poly35_ch3_q_o_net;
  q_fofb_o <= q_fofb_o_net;
  q_monit_o <= q_monit_o_net;
  q_tbt_o <= q_tbt_o_net;
  sum_fofb_o <= sum_fofb_o_net;
  sum_monit_o <= sum_monit_o_net;
  sum_tbt_o <= sum_tbt_o_net;
  tbt_amp_ch0_o <= tbt_amp_ch0_o_net;
  tbt_amp_ch1_o <= tbt_amp_ch1_o_net;
  tbt_amp_ch2_o <= tbt_amp_ch2_o_net;
  tbt_amp_ch3_o <= tbt_amp_ch3_o_net;
  x_fofb_o <= x_fofb_o_net;
  x_monit_o <= x_monit_o_net;
  x_tbt_o <= x_tbt_o_net;
  y_fofb_o <= y_fofb_o_net;
  y_monit_o <= y_monit_o_net;
  y_tbt_o <= y_tbt_o_net;

  channel0_fofb_3577a252e5: entity work.channel0_fofb_entity_3577a252e5
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      mix_i_in => mix_ch0_i_o_net,
      mix_q_in => mix_ch0_q_o_net,
      amp_f => fofb_amp_ch0_o_net,
      cic_fofb_i_fpga_out => cic_fofb_ch0_i_o_net,
      cic_fofb_q_fpga_out => cic_fofb_ch0_q_o_net,
      valid_f => register6_q_net_x4
    );

  channel0_tbt_b3ebb9eccb: entity work.channel0_tbt_entity_b3ebb9eccb
    port map (
      adc_ch0_i => adc_ch0_i_net_x2,
      ce_1 => ce_1_sg_x48,
      ce_35 => ce_35_sg_x13,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_35 => clk_35_sg_x13,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x11,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x11,
      dds_valid_in => dds_m_axis_data_tvalid_net_x11,
      amp_f => tbt_amp_ch0_o_net,
      bpf_adc_fpga_out => bpf_ch0_o_net,
      decim_35_i_fpga_out => poly35_ch0_i_o_net,
      decim_35_q_fpga_out => poly35_ch0_q_o_net,
      mix_i => mix_ch0_i_o_net,
      mix_q => mix_ch0_q_o_net,
      valid_f => register6_q_net_x5
    );

  channel1_fofb_8f5127405d: entity work.channel0_fofb_entity_3577a252e5
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      mix_i_in => mix_ch1_i_o_net,
      mix_q_in => mix_ch1_q_o_net,
      amp_f => fofb_amp_ch1_o_net,
      cic_fofb_i_fpga_out => cic_fofb_ch1_i_o_net,
      cic_fofb_q_fpga_out => cic_fofb_ch1_q_o_net,
      valid_f => register6_q_net_x6
    );

  channel1_tbt_8d468f1125: entity work.channel1_tbt_entity_8d468f1125
    port map (
      adc_ch1_i => adc_ch1_i_net_x2,
      ce_1 => ce_1_sg_x48,
      ce_35 => ce_35_sg_x13,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_35 => clk_35_sg_x13,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x11,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x11,
      dds_valid_in => dds_m_axis_data_tvalid_net_x11,
      amp_f => tbt_amp_ch1_o_net,
      bpf_adc_fpga_out => bpf_ch1_o_net,
      decim_35_i_fpga_out => poly35_ch1_i_o_net,
      decim_35_q_fpga_out => poly35_ch1_q_o_net,
      mix_i => mix_ch1_i_o_net,
      mix_q => mix_ch1_q_o_net,
      valid_f => register6_q_net_x7
    );

  channel2_fofb_c122b5720b: entity work.channel0_fofb_entity_3577a252e5
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      mix_i_in => mix_ch2_i_o_net,
      mix_q_in => mix_ch2_q_o_net,
      amp_f => fofb_amp_ch2_o_net,
      cic_fofb_i_fpga_out => cic_fofb_ch2_i_o_net,
      cic_fofb_q_fpga_out => cic_fofb_ch2_q_o_net,
      valid_f => register6_q_net_x8
    );

  channel2_tbt_c5e2abdcfa: entity work.channel2_tbt_entity_c5e2abdcfa
    port map (
      adc_ch2_i => adc_ch2_i_net_x2,
      ce_1 => ce_1_sg_x48,
      ce_35 => ce_35_sg_x13,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_35 => clk_35_sg_x13,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x11,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x11,
      dds_valid_in => dds_m_axis_data_tvalid_net_x11,
      amp_f => tbt_amp_ch2_o_net,
      bpf_adc_fpga_out => bpf_ch2_o_net,
      decim_35_i_fpga_out => poly35_ch2_i_o_net,
      decim_35_q_fpga_out => poly35_ch2_q_o_net,
      mix_i => mix_ch2_i_o_net,
      mix_q => mix_ch2_q_o_net,
      valid_f => register6_q_net_x9
    );

  channel3_fofb_79576133ce: entity work.channel0_fofb_entity_3577a252e5
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      mix_i_in => mix_ch3_i_o_net,
      mix_q_in => mix_ch3_q_o_net,
      amp_f => fofb_amp_ch3_o_net,
      cic_fofb_i_fpga_out => cic_fofb_ch3_i_o_net,
      cic_fofb_q_fpga_out => cic_fofb_ch3_q_o_net,
      valid_f => register6_q_net_x10
    );

  channel3_tbt_63129db436: entity work.channel3_tbt_entity_63129db436
    port map (
      adc_ch3_i => adc_ch3_i_net_x2,
      ce_1 => ce_1_sg_x48,
      ce_35 => ce_35_sg_x13,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x48,
      clk_35 => clk_35_sg_x13,
      dds_cosine_in => dds_m_axis_data_tdata_cosine_net_x11,
      dds_msine_in => dds_m_axis_data_tdata_sine_net_x11,
      dds_valid_in => dds_m_axis_data_tvalid_net_x11,
      amp_f => tbt_amp_ch3_o_net,
      bpf_adc_fpga_out => bpf_ch3_o_net,
      decim_35_i_fpga_out => poly35_ch3_i_o_net,
      decim_35_q_fpga_out => poly35_ch3_q_o_net,
      mix_i => mix_ch3_i_o_net,
      mix_q => mix_ch3_q_o_net,
      valid_f => register6_q_net_x11
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  dds: entity work.xldds_compiler_b7bbc719459e4bb4074716a9175f7d86
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      m_axis_data_tready => constant3_op_net,
      m_axis_data_tdata_cosine => dds_m_axis_data_tdata_cosine_net_x11,
      m_axis_data_tdata_sine => dds_m_axis_data_tdata_sine_net_x11,
      m_axis_data_tvalid => dds_m_axis_data_tvalid_net_x11
    );

  decim_q_monit_d3ca57d66c: entity work.decim_q_monit_entity_d3ca57d66c
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_11130000 => ce_11130000_sg_x4,
      ce_2782500 => ce_2782500_sg_x4,
      ce_5565000 => ce_5565000_sg_x4,
      ce_logic_1113 => ce_logic_1113_sg_x4,
      ce_logic_2782500 => ce_logic_2782500_sg_x4,
      ce_logic_5565000 => ce_logic_5565000_sg_x4,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      clk_11130000 => clk_11130000_sg_x4,
      clk_2782500 => clk_2782500_sg_x4,
      clk_5565000 => clk_5565000_sg_x4,
      data_in => down_sample2_q_net_x0,
      monit_out => q_monit_o_net
    );

  decim_sum_monit_1ee5debdc8: entity work.decim_sum_monit_entity_1ee5debdc8
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_11130000 => ce_11130000_sg_x4,
      ce_2782500 => ce_2782500_sg_x4,
      ce_5565000 => ce_5565000_sg_x4,
      ce_logic_1113 => ce_logic_1113_sg_x4,
      ce_logic_2782500 => ce_logic_2782500_sg_x4,
      ce_logic_5565000 => ce_logic_5565000_sg_x4,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      clk_11130000 => clk_11130000_sg_x4,
      clk_2782500 => clk_2782500_sg_x4,
      clk_5565000 => clk_5565000_sg_x4,
      data_in => down_sample3_q_net_x0,
      monit_out => sum_monit_o_net
    );

  decim_x_monit_75f6043a5c: entity work.decim_q_monit_entity_d3ca57d66c
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_11130000 => ce_11130000_sg_x4,
      ce_2782500 => ce_2782500_sg_x4,
      ce_5565000 => ce_5565000_sg_x4,
      ce_logic_1113 => ce_logic_1113_sg_x4,
      ce_logic_2782500 => ce_logic_2782500_sg_x4,
      ce_logic_5565000 => ce_logic_5565000_sg_x4,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      clk_11130000 => clk_11130000_sg_x4,
      clk_2782500 => clk_2782500_sg_x4,
      clk_5565000 => clk_5565000_sg_x4,
      data_in => down_sample_q_net_x0,
      monit_out => x_monit_o_net
    );

  decim_y_monit_902fe6e273: entity work.decim_q_monit_entity_d3ca57d66c
    port map (
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      ce_11130000 => ce_11130000_sg_x4,
      ce_2782500 => ce_2782500_sg_x4,
      ce_5565000 => ce_5565000_sg_x4,
      ce_logic_1113 => ce_logic_1113_sg_x4,
      ce_logic_2782500 => ce_logic_2782500_sg_x4,
      ce_logic_5565000 => ce_logic_5565000_sg_x4,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      clk_11130000 => clk_11130000_sg_x4,
      clk_2782500 => clk_2782500_sg_x4,
      clk_5565000 => clk_5565000_sg_x4,
      data_in => down_sample1_q_net_x0,
      monit_out => y_monit_o_net
    );

  delta_sigma_fofb_ee61e649ea: entity work.delta_sigma_fofb_entity_ee61e649ea
    port map (
      a => fofb_amp_ch0_o_net,
      avalid => register6_q_net_x4,
      b => fofb_amp_ch1_o_net,
      bvalid => register6_q_net_x6,
      c => fofb_amp_ch2_o_net,
      ce_1 => ce_1_sg_x48,
      ce_1113 => ce_1113_sg_x17,
      clk_1 => clk_1_sg_x48,
      clk_1113 => clk_1113_sg_x17,
      cvalid => register6_q_net_x8,
      d => fofb_amp_ch3_o_net,
      delta_sigma_thres => del_sig_div_fofb_thres_i_net,
      dvalid => register6_q_net_x10,
      q => q_fofb_o_net,
      sum_x0 => sum_fofb_o_net,
      x => x_fofb_o_net,
      y => y_fofb_o_net
    );

  delta_sigma_tbt_bbfa8a8a69: entity work.delta_sigma_tbt_entity_bbfa8a8a69
    port map (
      a => tbt_amp_ch0_o_net,
      avalid => register6_q_net_x5,
      b => tbt_amp_ch1_o_net,
      bvalid => register6_q_net_x7,
      c => tbt_amp_ch2_o_net,
      ce_1 => ce_1_sg_x48,
      ce_35 => ce_35_sg_x13,
      clk_1 => clk_1_sg_x48,
      clk_35 => clk_35_sg_x13,
      cvalid => register6_q_net_x9,
      d => tbt_amp_ch3_o_net,
      delta_sigma_thres => del_sig_div_tbt_thres_i_net,
      dvalid => register6_q_net_x11,
      q => q_tbt_o_net,
      sum_x0 => sum_tbt_o_net,
      x => x_tbt_o_net,
      y => y_tbt_o_net
    );

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 23,
      d_width => 24,
      ds_ratio => 1113,
      latency => 1,
      phase => 1112,
      q_arith => xlSigned,
      q_bin_pt => 23,
      q_width => 24
    )
    port map (
      d => x_fofb_o_net,
      dest_ce => ce_1113_sg_x17,
      dest_clk => clk_1113_sg_x17,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 23,
      d_width => 24,
      ds_ratio => 1113,
      latency => 1,
      phase => 1112,
      q_arith => xlSigned,
      q_bin_pt => 23,
      q_width => 24
    )
    port map (
      d => y_fofb_o_net,
      dest_ce => ce_1113_sg_x17,
      dest_clk => clk_1113_sg_x17,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 23,
      d_width => 24,
      ds_ratio => 1113,
      latency => 1,
      phase => 1112,
      q_arith => xlSigned,
      q_bin_pt => 23,
      q_width => 24
    )
    port map (
      d => q_fofb_o_net,
      dest_ce => ce_1113_sg_x17,
      dest_clk => clk_1113_sg_x17,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  down_sample3: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 20,
      d_width => 24,
      ds_ratio => 1113,
      latency => 1,
      phase => 1112,
      q_arith => xlSigned,
      q_bin_pt => 20,
      q_width => 24
    )
    port map (
      d => sum_fofb_o_net,
      dest_ce => ce_1113_sg_x17,
      dest_clk => clk_1113_sg_x17,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample3_q_net_x0
    );

end structural;
