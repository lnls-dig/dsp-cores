-------------------------------------------------------------------------------
-- Title      : Generic Multiplier
-- Project    :
-------------------------------------------------------------------------------
-- File       : generic_multiplier.vhd
-- Author     : aylons  <aylons@LNLS190>
-- Company    :
-- Created    : 2014-02-25
-- Last update: 2015-10-15
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: A multiplier where each input and output widths are determined
-- by generics. The inputs may be both unsigned, one signed or both signed, and
-- the ouput always have only one sign bit + MSBs.
-------------------------------------------------------------------------------
-- Copyright (c) 2014
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-02-25  1.0      aylons  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

-------------------------------------------------------------------------------

entity generic_multiplier is

  generic (
    g_a_width : natural := 16;          -- width for each input.
    g_b_width : natural := 16;

    g_signed : boolean := true;  -- signed or unsigned multiplication? Signed
    -- multiplication will have only one sign bit
    -- at the output

    g_p_width : natural := 16;          -- width for output. Must be less than
    -- g_a_width + g_b_width if unsigned,
    -- g_a_width+g_b_width-1 if signed.

    g_levels : natural := 7);           -- Just multiplier pipeline. Total
                                        -- delay is levels +2

  port (
    a_i     : in  std_logic_vector(g_a_width-1 downto 0);
    b_i     : in  std_logic_vector(g_b_width-1 downto 0);
    valid_i : in  std_logic;
    p_o     : out std_logic_vector(g_p_width-1 downto 0);
    valid_o : out std_logic;
    ce_i    : in  std_logic;
    clk_i   : in  std_logic;
    reset_i : in  std_logic);

  attribute mult_style                       : string;
  attribute mult_style of generic_multiplier : entity is "pipe_block";

end entity generic_multiplier;

-------------------------------------------------------------------------------

architecture behavioural of generic_multiplier is
  constant c_product_width : natural := g_a_width + g_b_width;

  type pipe is array(g_levels-1 downto 0) of std_logic_vector(c_product_width-1 downto 0);
  type pipe_valid is array(g_levels-1 downto 0) of std_logic;

  signal a       : std_logic_vector(g_a_width-1 downto 0) := (others => '0');
  signal b       : std_logic_vector(g_b_width-1 downto 0) := (others => '0');
  signal valid_in : std_logic                             := '0';
  signal product : pipe                                   := (others => (others => '0'));
  signal product_full : std_logic_vector(c_product_width-1 downto 0) := (others => '0');
  signal valid   : pipe_valid                             := (others => '0');
begin  -- architecture str

  -----------------------------------------------------------------------------
  -- Component instantiations
  -----------------------------------------------------------------------------

  -- Last stage of multiplication pipeline
  product_full <= product(g_levels-1);

  multiplication : process(clk_i)

  begin
    if rising_edge(clk_i) then

      if reset_i = '1' then
        p_o <= (others => '0');
        valid_o <= '0';

      elsif ce_i = '1' then

        -- Instantiate a register before multiplier to improve speed
        a <= a_i;
        b <= b_i;
        valid_in <= valid_i;

        -- If both are signed, there are two signals. Drop the redundancy.
        if g_signed = true then
          product(0) <= std_logic_vector(signed(a) * signed(b));
          valid(0) <= valid_in;
          for n in 1 to g_levels-1 loop
            product(n) <= product(n-1);
            valid(n) <= valid(n-1);
          end loop;

          if g_p_width < c_product_width then
            p_o <= product_full(c_product_width-2 downto c_product_width - g_p_width - 1);
            -- Keep "valid_o" grouped with "p_o" so we don't forget to keep them synchronized
            valid_o <= valid(g_levels-1);
          else
            p_o <= std_logic_vector(resize(signed(product_full), g_p_width));
            -- Keep "valid_o" grouped with "p_o" so we don't forget to keep them synchronized
            valid_o <= valid(g_levels-1);
          end if;


        else
          product(0) <= std_logic_vector(unsigned(a) * unsigned(b));
          valid(0) <= valid_in;

          for n in 1 to g_levels-1 loop
            product(n) <= product(n-1);
            valid(n) <= valid(n-1);
          end loop;

          if g_p_width < c_product_width then
            p_o <= product_full(c_product_width-1 downto c_product_width - g_p_width);
            -- Keep "valid_o" grouped with "p_o" so we don't forget to keep them synchronized
            valid_o <= valid(g_levels-1);
          else
            p_o <= std_logic_vector(resize(signed(product_full), g_p_width));
            -- Keep "valid_o" grouped with "p_o" so we don't forget to keep them synchronized
            valid_o <= valid(g_levels-1);
          end if;

        end if;

      end if;  -- reset
    end if;  -- clk
  end process multiplication;

end architecture behavioural;

-------------------------------------------------------------------------------
