--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_293aa5f110d040c2.vhd when simulating
-- the core, addsb_11_0_293aa5f110d040c2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_293aa5f110d040c2 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(24 DOWNTO 0)
  );
END addsb_11_0_293aa5f110d040c2;

ARCHITECTURE addsb_11_0_293aa5f110d040c2_a OF addsb_11_0_293aa5f110d040c2 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_293aa5f110d040c2
  PORT (
    a : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(24 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_293aa5f110d040c2 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 25,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000000000000000",
      c_b_width => 25,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 25,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_293aa5f110d040c2
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_293aa5f110d040c2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_3537d66a2361cd1e.vhd when simulating
-- the core, addsb_11_0_3537d66a2361cd1e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_3537d66a2361cd1e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END addsb_11_0_3537d66a2361cd1e;

ARCHITECTURE addsb_11_0_3537d66a2361cd1e_a OF addsb_11_0_3537d66a2361cd1e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_3537d66a2361cd1e
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_3537d66a2361cd1e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 26,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000000000",
      c_b_width => 26,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 26,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_3537d66a2361cd1e
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_3537d66a2361cd1e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_44053abf11139d96.vhd when simulating
-- the core, addsb_11_0_44053abf11139d96. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_44053abf11139d96 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END addsb_11_0_44053abf11139d96;

ARCHITECTURE addsb_11_0_44053abf11139d96_a OF addsb_11_0_44053abf11139d96 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_44053abf11139d96
  PORT (
    a : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(25 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(25 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_44053abf11139d96 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 26,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "00000000000000000000000000",
      c_b_width => 26,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 26,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_44053abf11139d96
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_44053abf11139d96_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cc_cmplr_v3_0_964aa42461b15ac2.vhd when simulating
-- the core, cc_cmplr_v3_0_964aa42461b15ac2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cc_cmplr_v3_0_964aa42461b15ac2 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END cc_cmplr_v3_0_964aa42461b15ac2;

ARCHITECTURE cc_cmplr_v3_0_964aa42461b15ac2_a OF cc_cmplr_v3_0_964aa42461b15ac2 IS
-- synthesis translate_off
COMPONENT wrapped_cc_cmplr_v3_0_964aa42461b15ac2
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cc_cmplr_v3_0_964aa42461b15ac2 USE ENTITY XilinxCoreLib.cic_compiler_v3_0(behavioral)
    GENERIC MAP (
      c_c1 => 58,
      c_c2 => 58,
      c_c3 => 58,
      c_c4 => 0,
      c_c5 => 0,
      c_c6 => 0,
      c_clk_freq => 2,
      c_component_name => "cc_cmplr_v3_0_964aa42461b15ac2",
      c_diff_delay => 2,
      c_family => "artix7",
      c_filter_type => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_dout_tready => 0,
      c_has_rounding => 0,
      c_i1 => 58,
      c_i2 => 58,
      c_i3 => 58,
      c_i4 => 0,
      c_i5 => 0,
      c_i6 => 0,
      c_input_width => 24,
      c_m_axis_data_tdata_width => 64,
      c_m_axis_data_tuser_width => 16,
      c_max_rate => 1120,
      c_min_rate => 1120,
      c_num_channels => 2,
      c_num_stages => 3,
      c_output_width => 58,
      c_rate => 1120,
      c_rate_type => 0,
      c_s_axis_config_tdata_width => 1,
      c_s_axis_data_tdata_width => 24,
      c_sample_freq => 1,
      c_use_dsp => 1,
      c_use_streaming_interface => 1,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cc_cmplr_v3_0_964aa42461b15ac2
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tdata => s_axis_data_tdata,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tlast => s_axis_data_tlast,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tlast => m_axis_data_tlast,
    event_tlast_unexpected => event_tlast_unexpected,
    event_tlast_missing => event_tlast_missing
  );
-- synthesis translate_on

END cc_cmplr_v3_0_964aa42461b15ac2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cc_cmplr_v3_0_e58a4eb9f6488d2d.vhd when simulating
-- the core, cc_cmplr_v3_0_e58a4eb9f6488d2d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cc_cmplr_v3_0_e58a4eb9f6488d2d IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END cc_cmplr_v3_0_e58a4eb9f6488d2d;

ARCHITECTURE cc_cmplr_v3_0_e58a4eb9f6488d2d_a OF cc_cmplr_v3_0_e58a4eb9f6488d2d IS
-- synthesis translate_off
COMPONENT wrapped_cc_cmplr_v3_0_e58a4eb9f6488d2d
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cc_cmplr_v3_0_e58a4eb9f6488d2d USE ENTITY XilinxCoreLib.cic_compiler_v3_0(behavioral)
    GENERIC MAP (
      c_c1 => 61,
      c_c2 => 61,
      c_c3 => 61,
      c_c4 => 0,
      c_c5 => 0,
      c_c6 => 0,
      c_clk_freq => 2240,
      c_component_name => "cc_cmplr_v3_0_e58a4eb9f6488d2d",
      c_diff_delay => 2,
      c_family => "artix7",
      c_filter_type => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_dout_tready => 0,
      c_has_rounding => 0,
      c_i1 => 61,
      c_i2 => 61,
      c_i3 => 61,
      c_i4 => 0,
      c_i5 => 0,
      c_i6 => 0,
      c_input_width => 24,
      c_m_axis_data_tdata_width => 64,
      c_m_axis_data_tuser_width => 16,
      c_max_rate => 2500,
      c_min_rate => 2500,
      c_num_channels => 4,
      c_num_stages => 3,
      c_output_width => 61,
      c_rate => 2500,
      c_rate_type => 0,
      c_s_axis_config_tdata_width => 1,
      c_s_axis_data_tdata_width => 24,
      c_sample_freq => 1,
      c_use_dsp => 1,
      c_use_streaming_interface => 1,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cc_cmplr_v3_0_e58a4eb9f6488d2d
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tdata => s_axis_data_tdata,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tlast => s_axis_data_tlast,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tlast => m_axis_data_tlast,
    event_tlast_unexpected => event_tlast_unexpected,
    event_tlast_missing => event_tlast_missing
  );
-- synthesis translate_on

END cc_cmplr_v3_0_e58a4eb9f6488d2d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cmpy_v5_0_02d02e0a23eb9773.vhd when simulating
-- the core, cmpy_v5_0_02d02e0a23eb9773. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cmpy_v5_0_02d02e0a23eb9773 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_a_tvalid : IN STD_LOGIC;
    s_axis_a_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    s_axis_b_tvalid : IN STD_LOGIC;
    s_axis_b_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_b_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END cmpy_v5_0_02d02e0a23eb9773;

ARCHITECTURE cmpy_v5_0_02d02e0a23eb9773_a OF cmpy_v5_0_02d02e0a23eb9773 IS
-- synthesis translate_off
COMPONENT wrapped_cmpy_v5_0_02d02e0a23eb9773
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_a_tvalid : IN STD_LOGIC;
    s_axis_a_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    s_axis_b_tvalid : IN STD_LOGIC;
    s_axis_b_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_b_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cmpy_v5_0_02d02e0a23eb9773 USE ENTITY XilinxCoreLib.cmpy_v5_0(behavioral)
    GENERIC MAP (
      c_a_width => 24,
      c_b_width => 24,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_s_axis_a_tlast => 0,
      c_has_s_axis_a_tuser => 0,
      c_has_s_axis_b_tlast => 0,
      c_has_s_axis_b_tuser => 1,
      c_has_s_axis_ctrl_tlast => 0,
      c_has_s_axis_ctrl_tuser => 0,
      c_latency => 6,
      c_m_axis_dout_tdata_width => 48,
      c_m_axis_dout_tuser_width => 1,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_width => 24,
      c_s_axis_a_tdata_width => 48,
      c_s_axis_a_tuser_width => 1,
      c_s_axis_b_tdata_width => 48,
      c_s_axis_b_tuser_width => 1,
      c_s_axis_ctrl_tdata_width => 8,
      c_s_axis_ctrl_tuser_width => 1,
      c_throttle_scheme => 3,
      c_tlast_resolution => 0,
      c_verbosity => 0,
      c_xdevice => "xc7a200t",
      c_xdevicefamily => "artix7",
      has_negate => 0,
      round => 0,
      single_output => 0,
      use_dsp_cascades => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cmpy_v5_0_02d02e0a23eb9773
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_a_tvalid => s_axis_a_tvalid,
    s_axis_a_tdata => s_axis_a_tdata,
    s_axis_b_tvalid => s_axis_b_tvalid,
    s_axis_b_tuser => s_axis_b_tuser,
    s_axis_b_tdata => s_axis_b_tdata,
    m_axis_dout_tvalid => m_axis_dout_tvalid,
    m_axis_dout_tuser => m_axis_dout_tuser,
    m_axis_dout_tdata => m_axis_dout_tdata
  );
-- synthesis translate_on

END cmpy_v5_0_02d02e0a23eb9773_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_eb46eda57512a5a4.vhd when simulating
-- the core, cntr_11_0_eb46eda57512a5a4. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_eb46eda57512a5a4 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END cntr_11_0_eb46eda57512a5a4;

ARCHITECTURE cntr_11_0_eb46eda57512a5a4_a OF cntr_11_0_eb46eda57512a5a4 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_eb46eda57512a5a4
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_eb46eda57512a5a4 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 2,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_eb46eda57512a5a4
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_eb46eda57512a5a4_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file crdc_v5_0_3d2446e74ce31176.vhd when simulating
-- the core, crdc_v5_0_3d2446e74ce31176. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY crdc_v5_0_3d2446e74ce31176 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_cartesian_tvalid : IN STD_LOGIC;
    s_axis_cartesian_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_cartesian_tdata : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END crdc_v5_0_3d2446e74ce31176;

ARCHITECTURE crdc_v5_0_3d2446e74ce31176_a OF crdc_v5_0_3d2446e74ce31176 IS
-- synthesis translate_off
COMPONENT wrapped_crdc_v5_0_3d2446e74ce31176
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_cartesian_tvalid : IN STD_LOGIC;
    s_axis_cartesian_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_cartesian_tdata : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    m_axis_dout_tvalid : OUT STD_LOGIC;
    m_axis_dout_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_dout_tdata : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_crdc_v5_0_3d2446e74ce31176 USE ENTITY XilinxCoreLib.cordic_v5_0(behavioral)
    GENERIC MAP (
      c_architecture => 2,
      c_coarse_rotate => 1,
      c_cordic_function => 1,
      c_data_format => 0,
      c_has_aclk => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_s_axis_cartesian => 1,
      c_has_s_axis_cartesian_tlast => 0,
      c_has_s_axis_cartesian_tuser => 1,
      c_has_s_axis_phase => 0,
      c_has_s_axis_phase_tlast => 0,
      c_has_s_axis_phase_tuser => 0,
      c_input_width => 25,
      c_iterations => 0,
      c_m_axis_dout_tdata_width => 48,
      c_m_axis_dout_tuser_width => 1,
      c_output_width => 24,
      c_phase_format => 0,
      c_pipeline_mode => -1,
      c_precision => 0,
      c_round_mode => 3,
      c_s_axis_cartesian_tdata_width => 64,
      c_s_axis_cartesian_tuser_width => 1,
      c_s_axis_phase_tdata_width => 32,
      c_s_axis_phase_tuser_width => 1,
      c_scale_comp => 3,
      c_throttle_scheme => 3,
      c_tlast_resolution => 0,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_crdc_v5_0_3d2446e74ce31176
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_cartesian_tvalid => s_axis_cartesian_tvalid,
    s_axis_cartesian_tuser => s_axis_cartesian_tuser,
    s_axis_cartesian_tdata => s_axis_cartesian_tdata,
    m_axis_dout_tvalid => m_axis_dout_tvalid,
    m_axis_dout_tuser => m_axis_dout_tuser,
    m_axis_dout_tdata => m_axis_dout_tdata
  );
-- synthesis translate_on

END crdc_v5_0_3d2446e74ce31176_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.87xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v4_0_dc31160d1288a80d.vhd
-- /___/   /\     Timestamp: Mon Sep 30 17:15:10 2013
-- \   \  /  \
--  \___\/\___\
--
-- Command	: -w -sim -ofmt vhdl C:/TEMP/sysgentmp-lucas.russo/cg_wk/c66822aecbec157bb/tmp/_cg/dv_gn_v4_0_dc31160d1288a80d.ngc C:/TEMP/sysgentmp-lucas.russo/cg_wk/c66822aecbec157bb/tmp/_cg/dv_gn_v4_0_dc31160d1288a80d.vhd
-- Device	: 7a200tffg1156-1
-- Input file	: C:/TEMP/sysgentmp-lucas.russo/cg_wk/c66822aecbec157bb/tmp/_cg/dv_gn_v4_0_dc31160d1288a80d.ngc
-- Output file	: C:/TEMP/sysgentmp-lucas.russo/cg_wk/c66822aecbec157bb/tmp/_cg/dv_gn_v4_0_dc31160d1288a80d.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v4_0_dc31160d1288a80d
-- Xilinx	: c:\xilinx\13.4\ise_ds\ise\
--
-- Purpose:
--     This VHDL netlist is a verification model and uses simulation
--     primitives which may not represent the true implementation of the
--     device, however the netlist is functionally correct and should not
--     be modified. This file cannot be synthesized and should only be used
--     with supported simulation tools.
--
-- Reference:
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v4_0_dc31160d1288a80d is
  port (
    aclk : in STD_LOGIC := 'X';
    aclken : in STD_LOGIC := 'X';
    s_axis_divisor_tvalid : in STD_LOGIC := 'X';
    s_axis_dividend_tvalid : in STD_LOGIC := 'X';
    s_axis_divisor_tready : out STD_LOGIC;
    s_axis_dividend_tready : out STD_LOGIC;
    m_axis_dout_tvalid : out STD_LOGIC;
    s_axis_divisor_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    s_axis_dividend_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    m_axis_dout_tdata : out STD_LOGIC_VECTOR ( 55 downto 0 )
  );
end dv_gn_v4_0_dc31160d1288a80d;

architecture STRUCTURE of dv_gn_v4_0_dc31160d1288a80d is
  signal NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_valid_access_in : STD_LOGIC;
  signal U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_56_110 : STD_LOGIC;
  signal U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_quot_det : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_sync_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_sync_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_start_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_start_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_3_374 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_4_375 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_3_376 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_4_377 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_3_378 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_4_379 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_pre_a : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_rfd : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_27_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_28_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_50_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_49_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_40_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_41_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_42_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_43_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_44_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_45_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_46_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_47_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_47_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_46_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_45_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_44_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_43_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_42_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_41_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_39_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_38_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_37_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_36_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_35_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_34_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_33_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_31_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_30_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_29_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_28_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_27_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_26_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_25_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_23_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_22_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_21_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_20_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_19_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_18_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_17_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_15_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_14_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_13_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_12_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_11_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_10_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_9_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_7_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_6_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_5_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_4_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_3_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_2_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_1_inv_not_gen_inv_thr_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_0_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_1_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_2_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_3_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_4_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_5_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_6_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_7_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_8_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_9_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_10_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_11_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_12_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_13_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_14_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_15_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_16_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_17_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_18_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_19_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_20_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_21_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_22_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_23_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_24_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_25_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_4_del_ce_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_3_del_ce_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_2_del_ce_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_0_del_ce_opt_has_pipe_first_q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_Mxor_quot_det_xo_0_1_2086 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_rt_2087 : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_rt_2088 : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_rt_2089 : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_rt_2090 : STD_LOGIC;

  signal N2 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0_2092 : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1_2093 : STD_LOGIC;

  signal U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0_2094 : STD_LOGIC;
  signal U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1_2095 : STD_LOGIC;
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0_2096 : STD_LOGIC;

  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1_2097 : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0_Q_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1_Q31_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0_Q_UNCONNECTED : STD_LOGIC;
  signal NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1_Q31_UNCONNECTED : STD_LOGIC;
  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0_Q_UNCONNECTED : STD_LOGIC;

  signal NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1_Q31_UNCONNECTED : STD_LOGIC;

  signal NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i : STD_LOGIC_VECTOR ( 25 downto 25 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 50 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53 : STD_LOGIC_VECTOR ( 1 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i : STD_LOGIC_VECTOR ( 25 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i : STD_LOGIC_VECTOR ( 25 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i : STD_LOGIC_VECTOR ( 25 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a : STD_LOGIC_VECTOR ( 24 downto 1 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i : STD_LOGIC_VECTOR ( 25 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a : STD_LOGIC_VECTOR ( 24 downto 1 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 1 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase : STD_LOGIC_VECTOR ( 2 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result : STD_LOGIC_VECTOR ( 2 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi : STD_LOGIC_VECTOR ( 50 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q : STD_LOGIC_VECTOR ( 50 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i : STD_LOGIC_VECTOR ( 25 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a : STD_LOGIC_VECTOR ( 25 downto 1 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy : STD_LOGIC_VECTOR ( 23 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i : STD_LOGIC_VECTOR ( 24 downto 0 );
  signal U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a : STD_LOGIC_VECTOR ( 23 downto 1 );
begin
  m_axis_dout_tdata(55) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(54) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(53) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(52) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(51) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(50) <=
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25);
  m_axis_dout_tdata(49) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(24);
  m_axis_dout_tdata(48) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(23);
  m_axis_dout_tdata(47) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(22);
  m_axis_dout_tdata(46) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(21);
  m_axis_dout_tdata(45) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(20);
  m_axis_dout_tdata(44) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(19);
  m_axis_dout_tdata(43) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(18);
  m_axis_dout_tdata(42) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(17);
  m_axis_dout_tdata(41) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(16);
  m_axis_dout_tdata(40) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(15);
  m_axis_dout_tdata(39) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(14);
  m_axis_dout_tdata(38) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(13);
  m_axis_dout_tdata(37) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(12);
  m_axis_dout_tdata(36) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(11);
  m_axis_dout_tdata(35) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(10);
  m_axis_dout_tdata(34) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(9);
  m_axis_dout_tdata(33) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(8);
  m_axis_dout_tdata(32) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(7);
  m_axis_dout_tdata(31) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(6);
  m_axis_dout_tdata(30) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(5);
  m_axis_dout_tdata(29) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(4);
  m_axis_dout_tdata(28) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(3);
  m_axis_dout_tdata(27) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(2);
  m_axis_dout_tdata(26) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(1);
  m_axis_dout_tdata(25) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(0);
  m_axis_dout_tdata(24) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(24);
  m_axis_dout_tdata(23) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(23);
  m_axis_dout_tdata(22) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(22);
  m_axis_dout_tdata(21) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(21);
  m_axis_dout_tdata(20) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(20);
  m_axis_dout_tdata(19) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(19);
  m_axis_dout_tdata(18) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(18);
  m_axis_dout_tdata(17) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(17);
  m_axis_dout_tdata(16) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(16);
  m_axis_dout_tdata(15) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(15);
  m_axis_dout_tdata(14) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(14);
  m_axis_dout_tdata(13) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(13);
  m_axis_dout_tdata(12) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(12);
  m_axis_dout_tdata(11) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(11);
  m_axis_dout_tdata(10) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(10);
  m_axis_dout_tdata(9) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(9);
  m_axis_dout_tdata(8) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(8);
  m_axis_dout_tdata(7) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(7);
  m_axis_dout_tdata(6) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(6);
  m_axis_dout_tdata(5) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(5);
  m_axis_dout_tdata(4) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(4);
  m_axis_dout_tdata(3) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(3);
  m_axis_dout_tdata(2) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(2);
  m_axis_dout_tdata(1) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(1);
  m_axis_dout_tdata(0) <=
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(0);
  s_axis_divisor_tready <=
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q;
  s_axis_dividend_tready <=
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q;
  XST_GND : GND
    port map (
      G =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_valid_access_in,
      Q => U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_start_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => s_axis_dividend_tdata(25),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_start_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_start_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => s_axis_divisor_tdata(25),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_start_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_sync_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_start_opt_has_pipe_first_q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_sync_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_sync_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_start_opt_has_pipe_first_q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_sync_opt_has_pipe_first_q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_25_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(24),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_24_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(23),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_24_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(23),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(24)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_23_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(22),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_23_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(22),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(23)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_22_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(21),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_22_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(21),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(22)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_21_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(20),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_21_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(20),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(21)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_20_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(19),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_20_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(19),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(20)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_19_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(18),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_19_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(18),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(19)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_18_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(17),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_18_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(17),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(18)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_17_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(16),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_17_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(16),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(17)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_16_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(15),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_16_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(15),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(16)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_15_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(14),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_15_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(14),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(15)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_14_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(13),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_14_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(13),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(14)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_13_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(12),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_13_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(12),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(13)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_12_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(11),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_12_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(11),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(12)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_11_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(10),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_11_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(10),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(11)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_10_Q :
XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(9)
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_10_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(9)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(10)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_9_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(8)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(9)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_9_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(8)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_8_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(7)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(8)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_8_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(7)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_7_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(6)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(7)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_7_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(6)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_6_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(5)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(6)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_6_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(5)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_5_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(4)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(5)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_5_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(4)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_4_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(3)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(4)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_4_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(3)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_3_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(2)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(3)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_3_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(2)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_2_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(1)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(2)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_2_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(1)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_1_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(0)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(1)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_1_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(0)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_xor_0_Q : XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_rt_2087,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      DI => s_axis_dividend_tdata(25),
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_rt_2087,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(25),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(24),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(23),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(22),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(21),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(20),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(19),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_s_i(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_25_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(24)
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_24_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(23)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(24)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_24_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(23)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_23_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(22)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(23)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_23_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(22)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_22_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(21)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(22)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_22_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(21)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_21_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(20)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(21)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_21_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(20)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_20_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(19)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(20)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_20_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(19)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_19_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(18)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(19)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_19_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(18)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_18_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(17)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(18)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_18_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(17)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_17_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(16)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(17)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_17_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(16)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_16_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(15)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(16)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_16_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(15)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_15_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(14)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(15)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_15_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(14)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_14_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(13)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(14)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_14_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(13)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_13_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(12)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(13)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_13_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(12)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_12_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(11)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(12)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_12_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(11)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_11_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(10)
,
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(11)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_11_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(10)
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_10_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(9),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(10)
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_10_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(9),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_9_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(8),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_9_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(8),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_8_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(7),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_8_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(7),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_7_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(6),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_7_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(6),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_6_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(5),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_6_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(5),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_5_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(4),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_5_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(4),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_4_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(3),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_4_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(3),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_3_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(2),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_3_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(2),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_2_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(1),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_2_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(1),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_1_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(0),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_1_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(0),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_xor_0_Q : XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_rt_2088,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      DI => s_axis_divisor_tdata(25),
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_rt_2088,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(25),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(24),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(23),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(22),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(21),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(20),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(19),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i_0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_s_i(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_dividend_sync_opt_has_pipe_first_q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_msb_divisor_sync_opt_has_pipe_first_q,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_3 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_3_374
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_4 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_4_375
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_2_f7 : MUXF7
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_4_375,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_16_3_374,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_3 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_3_376
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_4 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_4_377
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_2_f7 : MUXF7
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_4_377,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_8_3_376,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_3 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_19_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_18_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_20_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_3_378
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_4 : LUT6
    generic map(
      INIT => X"FD75B931EC64A820"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_23_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_22_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_24_Q
,
      I5 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_4_379
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_2_f7 : MUXF7
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_4_379,
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_numer_mux_0_3_378,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_1_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_1_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_2_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_1_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_2_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_3_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_2_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_3_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_4_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_3_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_4_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_5_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_4_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_5_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_6_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_5_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_6_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_7_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_6_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_7_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_9_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_9_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_10_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_9_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_10_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_11_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_10_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_11_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_12_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_11_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_12_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_13_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_12_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_13_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_14_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_13_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_14_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_15_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_14_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_15_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_17_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_17_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_18_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_17_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_18_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_19_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_18_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_19_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_20_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_19_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_20_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_21_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_20_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_21_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_22_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_21_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_22_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_23_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_22_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_23_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_25_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_25_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_26_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_25_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_26_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_27_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_26_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_27_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_28_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_27_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_28_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_29_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_28_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_29_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_30_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_29_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_30_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_31_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_30_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_31_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_33_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_33_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_34_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_33_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_34_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_35_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_34_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_35_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_36_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_35_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_36_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_37_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_36_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_37_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_38_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_37_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_38_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_39_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_38_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_39_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_41_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_41_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_42_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_41_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_42_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_43_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_42_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_43_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_44_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_43_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_44_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_45_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_44_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_45_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_46_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_45_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_46_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_47_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_46_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_47_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_49_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_49_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_50_inv_not_gen_inv_thr_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_49_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_50_inv_not_gen_inv_thr_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(2),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_rfd,
      Q =>
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_0_del_ce_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_pre_a,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_0_del_ce_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_0_del_ce_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_2_del_ce_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_2_del_ce_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_3_del_ce_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_2_del_ce_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_3_del_ce_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_4_del_ce_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_3_del_ce_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_4_del_ce_opt_has_pipe_first_q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(25),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(24),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(23),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(22),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(21),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(20),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(19),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(18),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(17),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(16),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(15),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(14),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(13),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(12),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(11),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(10),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(9),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(8),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(7),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(6),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(5),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(4),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(3),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(2),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(1),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_q_i(0),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(25),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(24),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(23),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(22),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(21),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(20),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(19),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(18),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(17),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(16),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(15),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(14),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(13),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(12),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(11),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(10),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(9),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(8),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(7),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(6),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(5),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(4),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(3),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(2),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(1),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_q_i(0),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_div_start_other_del_divisor_init_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_28_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_27_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_25_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_24_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_23_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_22_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_21_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_20_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_19_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_18_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_17_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_16_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_15_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_14_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_13_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_12_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_11_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_10_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_9_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_8_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_7_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_6_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_5_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_4_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_3_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_1_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_0_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carryxortop :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_2_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carryxor :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_25_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_24_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_23_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_22_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_21_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_20_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_19_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_18_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_17_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_16_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_15_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_14_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_13_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_12_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_11_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_10_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_9_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_8_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_7_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_6_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_5_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_4_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_3_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_2_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_carrychaingen_1_carrymux :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_25_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q
,
      O =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_gt_1_muxtop_carrymuxtop_O_UNCONNECTED

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_carryxor0 :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_i_need_mux_carrymux0 :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_0_Q
,
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_carry_simple_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_7_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_6_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_5_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_4_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_3_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_2_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_1_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_15_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_14_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_13_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_12_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_11_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_10_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_9_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_23_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_22_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_21_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_20_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_19_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_18_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_17_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_31_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_30_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_29_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_28_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_27_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_26_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_25_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_39_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_38_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_37_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_36_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_35_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_34_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_33_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_47 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_47_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_46 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_46_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_45 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_45_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_44 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_44_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_43 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_43_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_42 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_42_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_41 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_41_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_40 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_40_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_47_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_46_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_45_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_44_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_43_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_42_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_41_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_50 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_47_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(50)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_49 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_46_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(49)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_48 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_45_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(48)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_47 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_44_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(47)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_46 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_43_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(46)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_45 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_42_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(45)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_44 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_41_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(44)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_43 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_40_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(43)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_42 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_39_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(42)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_41 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_38_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(41)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_40 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_37_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(40)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_39 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_36_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(39)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_38 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_35_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(38)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_37 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_34_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(37)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_36 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_33_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(36)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_35 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_32_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(35)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_34 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_31_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(34)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_33 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_30_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(33)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_32 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_29_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(32)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_31 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_28_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(31)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_30 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_27_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(30)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_29 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_26_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(29)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_25_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(28)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_24_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(27)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_23_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_22_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_21_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_20_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_19_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_18_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_17_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_16_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_15_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_14_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_13_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_12_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_11_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_10_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_9_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_8_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_7_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_6_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_5_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_4_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_3_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_2_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_1_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_quot_gen_quot_reg_quot_out_opt_has_pipe_first_q_0_Q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_50_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_49_inv_not_gen_inv_thr_opt_has_pipe_first_q
,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q_0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_50 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(50),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(50)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_49 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(49),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(49)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_48 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(48),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(48)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_47 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(47),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(47)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_46 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(46),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(46)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_45 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(45),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(45)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_44 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(44),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(44)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_43 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(43),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(43)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_42 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(42),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(42)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_41 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(41),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(41)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_40 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(40),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(40)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_39 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(39),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(39)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_38 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(38),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(38)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_37 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(37),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(37)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_36 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(36),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(36)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_35 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(35),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(35)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_34 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(34),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(34)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_33 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(33),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(33)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_32 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(32),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(32)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_31 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(31),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(31)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_30 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(30),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(30)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_29 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(29),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(29)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_28 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(28),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(28)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_27 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(27),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(27)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_26 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(26),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_25 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(25),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_24 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(24),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_23 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(23),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_22 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(22),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_21 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(21),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_20 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(20),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_19 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(19),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_18 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(18),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_17 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(17),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_16 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(16),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_15 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(15),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_14 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(14),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_13 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(13),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_12 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(12),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_11 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(11),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_10 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(10),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_9 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(9),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_8 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(8),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_7 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(7),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_6 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(6),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_5 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(5),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_4 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(4),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_3 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(3),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_2 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(2),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_1 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(1),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q_0 :
FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(0),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_25_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(24),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_24_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(23),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_24_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(23),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_23_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(22),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_23_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(22),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_22_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(21),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_22_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(21),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_21_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(20),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_21_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(20),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_20_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(19),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_20_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(19),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_19_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(18),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_19_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(18),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_18_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(17),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_18_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(17),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_17_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(16),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_17_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(16),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_16_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(15),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_16_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(15),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_15_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(14),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_15_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(14),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_14_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(13),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_14_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(13),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_13_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(12),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_13_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(12),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_12_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(11),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_12_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(11),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_11_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(10),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_11_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(10),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_10_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(9),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_10_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(9),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_9_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(8),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_9_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(8),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_8_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(7),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_8_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(7),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_7_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(6),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_7_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(6),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_6_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(5),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_6_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(5),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_5_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(4),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_5_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(4),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_4_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(3),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_4_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(3),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_3_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(2),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_3_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(2),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_2_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(1),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_2_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(1),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_1_Q : XORCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(0),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_1_Q : MUXCY
    port map (
      CI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(0),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_xor_0_Q : XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_rt_2089,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_Q : MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_quot_det,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_rt_2089,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(25),
      Q =>
NlwRenamedSignal_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(24),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(23),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(22),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(21),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(20),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(19),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(18),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(17),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(16),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(15),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(14),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(13),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(12),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(11),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(10),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(9),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(8),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(7),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(6),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(5),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(4),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(3),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(2),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(1),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_s_i(0),
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_q_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_24_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(23),
      LI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_Mxor_quot_det_xo_0_1_2086,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_23_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(22),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(23),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_23_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(22),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(23),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_22_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(21),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(22),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_22_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(21),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(22),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_21_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(20),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(21),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_21_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(20),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(21),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_20_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(19),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(20),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_20_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(19),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(20),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_19_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(18),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(19),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_19_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(18),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(19),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_18_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(17),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(18),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_18_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(17),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(18),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_17_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(16),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(17),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_17_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(16),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(17),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_16_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(15),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(16),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_16_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(15),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(16),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_15_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(14),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(15),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_15_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(14),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(15),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_14_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(13),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(14),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_14_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(13),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(14),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_13_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(12),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(13),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_13_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(12),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(13),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_12_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(11),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(12),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_12_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(11),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(12),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_11_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(10),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(11),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_11_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(10),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(11),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_10_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(9),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(10),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_10_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(9),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(10),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_9_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(8),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_9_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(8),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(9),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_8_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(7),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_8_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(7),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(8),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_7_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(6),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_7_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(6),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(7),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_6_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(5),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_6_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(5),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(6),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_5_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(4),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_5_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(4),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(5),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_4_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(3),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_4_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(3),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(4),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_3_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(2),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_3_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(2),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(3),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_2_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(1),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_2_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(1),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(2),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_1_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(0),
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_1_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(0),
      DI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_xor_0_Q :
XORCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      LI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_rt_2090
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_Q :
MUXCY
    port map (
      CI =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      DI => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_quot_det,
      S =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_rt_2090
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(24),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(23),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(22),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(21),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(20),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(19),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(18),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(17),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(16),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(15),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(14),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(13),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(12),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(11),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(10),
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(9)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(8)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(7)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(6)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(5)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(4)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(3)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(2)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(1)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_s_i(0)
,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_q_i(0)
    );
  U0_i_synth_rdy_if1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => aclken,
      I1 => U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_56_110,
      O => m_axis_dout_tvalid
    );
  U0_i_synth_valid_access_in1 : LUT4
    generic map(
      INIT => X"8000"
    )
    port map (
      I0 => aclken,
      I1 =>
NlwRenamedSig_OI_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_rfd_timing_signed_d248_rfd_reg_del_rfd_opt_has_pipe_first_q
,
      I2 => s_axis_dividend_tvalid,
      I3 => s_axis_divisor_tvalid,
      O => U0_i_synth_valid_access_in
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_Mxor_quot_det_xo_0_1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_quot_det
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a28 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(1),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a31 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(10),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a41 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(11),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a51 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(12),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a61 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(13),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a71 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(14),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a81 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(15),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a91 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(16),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a101 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(17),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a111 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(18),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a121 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(19),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a131 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(2),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a141 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(20),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a151 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(21),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a161 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(22),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a171 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(23),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a181 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(24),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a211 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(3),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a221 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(4),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a231 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(5),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a241 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(6),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a251 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(7),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a261 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(8),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Mmux_simp_addp_a271 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_dividend_tdata(9),
      I1 => s_axis_dividend_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_simp_addp_a(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a28 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(1),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a31 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(10),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a41 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(11),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a51 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(12),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a61 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(13),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a71 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(14),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a81 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(15),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a91 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(16),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a101 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(17),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a111 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(18),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a121 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(19),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a131 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(2),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a141 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(20),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a151 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(21),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a161 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(22),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a171 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(23),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a181 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(24),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a211 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(3),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a221 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(4),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a231 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(5),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a241 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(6),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a251 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(7),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a261 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(8),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Mmux_simp_addp_a271 :
LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => s_axis_divisor_tdata(9),
      I1 => s_axis_divisor_tdata(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_simp_addp_a(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mcount_dclk_phase_xor_2_11 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(2),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_24_0_1 : LUT5
    generic map(
      INIT => X"11100100"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_1_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_numer_mux_ctrl_mux_cnt_del_opt_has_pipe_first_q_0_Q
,
      I3 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_1_Q
,
      I4 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_num_stages_numerator_gen_del_numer_opt_has_pipe_first_q_0_Q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_numer_mux_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mcount_dclk_phase_xor_1_11 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_pre_a_2_1 : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(2),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_pre_a
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_rfd_2_1 : LUT3
    generic map(
      INIT => X"08"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(2),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(1),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_rfd
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_4_del_ce_opt_has_pipe_first_q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_ce_sig_0_1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_0_del_ce_opt_has_pipe_first_q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_m
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_8_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_16_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_24_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_40_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_0_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_0_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_3_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_1_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_1_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_12_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_10_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_10_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_13_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_11_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_11_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_14_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_12_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_12_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_15_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_13_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_13_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_16_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_14_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_14_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_17_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_15_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_15_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_18_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_16_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_16_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_19_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_17_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_17_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_20_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_18_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_18_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_21_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_19_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_19_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_4_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_2_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_22_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_20_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_20_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_23_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_21_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_21_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_24_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_22_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_22_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_25_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_23_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_23_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_26_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_24_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_24_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_27_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_25_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_25_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_1 :
LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_28_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_26_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_5_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_3_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_3_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_6_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_4_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_4_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_7_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_5_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_5_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_8_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_6_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_6_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_9_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_7_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_7_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_10_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_8_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_8_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_1 :
LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_11_Q
,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_divisor_gen_divisor_dcother_del_divisor_opt_has_pipe_first_q_9_Q
,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_1_Q
,
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_48_adder_gen_no_reg_adsu_mod2_add1_no_pipelining_the_addsub_i_lut4_i_lut4_addsub_i_simple_model_halfsum_9_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_Mxor_quot_det_xo_0_11 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_Mxor_quot_det_xo_0_1_2086
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a21 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(26),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a131 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(27),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a27 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(2),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a221 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(28),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a131 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(3),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a231 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(29),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a201 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(4),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a241 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(30),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a211 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(5),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a251 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(31),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a221 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(6),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a261 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(32),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a231 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(7),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a271 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(33),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a241 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(8),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a281 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(34),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a251 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(9),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a31 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(35),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a261 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(10),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a41 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(36),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a31 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(11),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_29 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_29 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_210 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_210 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_210 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_13 : LUT3
    generic map(
      INIT => X"8F"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I1 => aclken,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_210 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_29 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_1_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_110 : LUT4
    generic map(
      INIT => X"087F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_110 : LUT4
    generic map(
      INIT => X"078F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_13 : LUT4
    generic map(
      INIT => X"087F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_13 : LUT4
    generic map(
      INIT => X"087F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_13 : LUT4
    generic map(
      INIT => X"087F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_110 : LUT4
    generic map(
      INIT => X"078F"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_26_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_26_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_0_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_211 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_211 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_221 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_221 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_221 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_221 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_211 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_25_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_25_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_28_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_201 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_201 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_211 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_211 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_211 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_211 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_201 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_24_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_24_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_27_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_191 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_191 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_201 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_201 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_201 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_201 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_191 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_23_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_23_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_26_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_181 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_181 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_191 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_191 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_191 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_191 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_181 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_22_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_22_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_25_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_171 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_171 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_181 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_181 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_181 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_181 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_171 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_21_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_21_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_24_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_161 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_161 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_171 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_171 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_171 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_171 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_161 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_20_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_20_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_23_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_151 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_151 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_161 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_161 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_161 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_161 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_151 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_19_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_19_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_22_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_141 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_141 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_151 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_151 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_151 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_151 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_141 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_18_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_18_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_21_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_131 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_131 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_141 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_141 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_141 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_141 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_131 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_17_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_17_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_20_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_121 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_121 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_121 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_121 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_121 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_121 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_121 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_16_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_16_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_19_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_111 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_111 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_111 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_111 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_111 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_111 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_111 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_15_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_15_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_18_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_101 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_101 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_101 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_101 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_101 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_101 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_101 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_14_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_14_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_17_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a51 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(37),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a41 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(12),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a61 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(38),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a51 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(13),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a71 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(39),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a61 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(14),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a81 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(40),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a71 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(15),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a91 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(41),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a81 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(16),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a101 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(42),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a91 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(17),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a111 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(43),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a101 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(18),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a121 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(44),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a111 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(19),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a141 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(45),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a121 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(20),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a151 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(46),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a141 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(21),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a161 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(47),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a151 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(22),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a171 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(48),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a161 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(23),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_91 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_91 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_91 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_91 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_91 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_91 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_91 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_13_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_13_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_16_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_81 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_81 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_81 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_81 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_81 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_81 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_81 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_12_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_12_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_15_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_71 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_71 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_71 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_71 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_71 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_71 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_71 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_11_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_11_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_14_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_61 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_61 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_61 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_61 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_61 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_61 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_61 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_10_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_10_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_13_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_51 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_51 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_51 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_51 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_51 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_51 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_51 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_9_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_9_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_12_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_41 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_41 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_41 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_41 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_41 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_41 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_41 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_8_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_8_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_11_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_31 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_31 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_31 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_31 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_31 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_31 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_31 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_7_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_7_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_10_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_281 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_281 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_291 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_291 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_291 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_291 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_281 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_6_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_6_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_9_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_271 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_271 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_281 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_281 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_281 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_281 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_271 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_5_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_5_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_8_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_261 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_261 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_271 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_271 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_271 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_271 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_261 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_4_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_4_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_7_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_251 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_251 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_261 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_261 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_261 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_261 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_251 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_3_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_3_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_6_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_241 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_241 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_251 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_251 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_251 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_251 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_241 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_2_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_2_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_5_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a181 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(49),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Mmux_simp_addp_a171 :
LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(24),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_simp_addp_a(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Mmux_simp_addp_a191 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(50),
      I1 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0),
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_simp_addp_a(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_231 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_231 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_241 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_241 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_241 : LUT4
    generic map(
      INIT => X"F780"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_241 : LUT3
    generic map(
      INIT => X"70"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_231 : LUT4
    generic map(
      INIT => X"F870"
    )
    port map (
      I0 => aclken,
      I1 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I2 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_1_Q,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_1_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_4_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_40_221 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_40_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_32_221 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_32_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_32_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_24_231 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_24_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_24_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_16_231 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_16_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_16_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_8_231 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_8_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_8_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_0_231 : LUT3
    generic map(
      INIT => X"2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_0_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_0_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mmux_pre_mux_o_48_221 : LUT4
    generic map(
      INIT => X"EA2A"
    )
    port map (
      I0 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_48_0_Q,
      I1 => aclken,
      I2 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_0_stage_zero_control_gen_ce_create_1_del_ce_opt_has_pipe_first_q
,
      I3 => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_adsu_o_40_0_Q,
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_pre_mux_o_48_3_Q
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => s_axis_dividend_tdata(0),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_dividend_twos_comp_Madd_s_i_cy_0_rt_2087
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => s_axis_divisor_tdata(0),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sgned_input_cmp_divisor_twos_comp_Madd_s_i_cy_0_rt_2088
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_rt : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(25),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_cmp_quot_twos_comp_Madd_s_i_cy_0_rt_2089
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_rt :
LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_reg_quot_out_reg_quot_opt_has_pipe_first_q(1),
      O =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_signed_output_remd_fract_cmp_remd_twos_comp_Madd_s_i_cy_0_rt_2090

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Mcount_dclk_phase_xor_0_11_INV_0 : INV
    port map (
      I => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_dclk_phase(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_Result(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_0_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(0),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(0)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_1_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(1),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(1)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_2_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(2),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(2)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_3_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(3),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(3)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_4_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(4),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(4)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_5_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(5),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(5)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_6_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(6),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(6)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_7_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(7),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(7)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_8_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(8),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(8)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_9_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(9),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(9)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_10_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(10),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(10)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_11_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(11),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(11)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_12_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(12),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(12)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_13_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(13),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(13)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_14_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(14),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(14)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_15_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(15),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(15)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_16_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(16),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(16)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_17_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(17),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(17)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_18_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(18),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(18)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_19_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(19),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(19)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_20_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(20),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(20)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_21_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(21),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(21)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_22_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(22),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(22)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_23_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(23),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(23)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_24_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(24),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(24)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_25_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(25),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(25)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_26_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(26),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(26)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_27_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(27),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(27)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_28_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(28),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(28)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_29_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(29),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(29)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_30_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(30),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(30)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_31_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(31),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(31)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_32_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(32),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(32)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_33_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(33),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(33)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_34_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(34),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(34)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_35_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(35),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(35)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_36_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(36),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(36)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_37_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(37),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(37)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_38_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(38),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(38)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_39_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(39),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(39)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_40_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(40),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(40)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_41_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(41),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(41)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_42_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(42),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(42)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_43_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(43),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(43)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_44_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(44),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(44)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_45_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(45),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(45)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_46_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(46),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(46)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_47_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(47),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(47)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_48_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(48),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(48)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_49_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(49),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(49)
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi_50_1_INV_0 : INV
    port map (
      I =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_final_sel_quot_sel_opt_has_pipe_first_q(50),
      O => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_qpi(50)
    );
  XST_VCC : VCC
    port map (
      P => N2
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0 :
SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q(0),
      CE => aclken,
      Q =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0_Q_UNCONNECTED
,
      Q31 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0_2092,
      A(4) => N2,
      A(3) => N2,
      A(2) => N2,
      A(1) => N2,
      A(0) => N2
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1 :
SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_0_2092,
      CE => aclken,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1_2093,
      Q31 =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1_Q31_UNCONNECTED
,
      A(4) => N2,
      A(3) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(2) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(1) => N2,
      A(0) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53_0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_0_1_2093,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(0)
    );
  U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nd_to_rdy_opt_has_pipe_first_q,
      CE => aclken,
      Q => NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0_Q_UNCONNECTED,
      Q31 => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0_2094,
      A(4) => N2,
      A(3) => N2,
      A(2) => N2,
      A(1) => N2,
      A(0) => N2
    );
  U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_0_2094,
      CE => aclken,
      Q => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1_2095,
      Q31 => NLW_U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1_Q31_UNCONNECTED,
      A(4) => N2,
      A(3) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(2) => N2,
      A(1) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(0) => N2
    );
  U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_56 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D => U0_i_synth_i_nd_to_rdy_Mshreg_opt_has_pipe_pipe_56_1_2095,
      Q => U0_i_synth_i_nd_to_rdy_opt_has_pipe_pipe_56_110
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0 :
SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_first_q(1),
      CE => aclken,
      Q =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0_Q_UNCONNECTED
,
      Q31 =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0_2096,
      A(4) => N2,
      A(3) => N2,
      A(2) => N2,
      A(1) => N2,
      A(0) => N2
    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1 :
SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_0_2096,
      CE => aclken,
      Q =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1_2097,
      Q31 =>
NLW_U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1_Q31_UNCONNECTED
,
      A(4) => N2,
      A(3) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(2) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q
,
      A(1) => N2,
      A(0) =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_divider_blk_div_loop_32_mux_div_clock_mux_sig_mux_adsu_opt_has_pipe_first_q_2_Q

    );
  U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53_1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => aclken,
      D =>
U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_Mshreg_opt_has_pipe_pipe_53_1_1_2097,
      Q => U0_i_synth_i_nonzero_fract_i_synth_i_algo_r2_nr_i_nonzero_fract_i_sdivider_I_SYNTH_MODEL_sign_pipeline_sign_pipe_opt_has_pipe_pipe_53(1)
    );

end STRUCTURE;

-- synthesis translate_on
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_15ffe94f3ff4129f.vhd when simulating
-- the core, fr_cmplr_v6_3_15ffe94f3ff4129f. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_15ffe94f3ff4129f IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END fr_cmplr_v6_3_15ffe94f3ff4129f;

ARCHITECTURE fr_cmplr_v6_3_15ffe94f3ff4129f_a OF fr_cmplr_v6_3_15ffe94f3ff4129f IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_15ffe94f3ff4129f
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_15ffe94f3ff4129f USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "41",
      c_accum_path_widths => "41",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_15ffe94f3ff4129f.mif",
      c_coef_file_lines => 42,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "1",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_15ffe94f3ff4129f",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 1,
      c_data_memtype => 1,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "24",
      c_data_width => 24,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 2800000,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 30,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 1,
      c_m_data_tdata_width => 32,
      c_m_data_tuser_width => 2,
      c_mem_arrangement => 1,
      c_num_channels => 4,
      c_num_filts => 1,
      c_num_madds => 1,
      c_num_reload_slots => 1,
      c_num_taps => 81,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "25",
      c_output_rate => 5600000,
      c_output_width => 25,
      c_oversampling_rate => 21,
      c_reload_tdata_width => 1,
      c_round_mode => 4,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 1,
      c_s_data_tdata_width => 24,
      c_s_data_tuser_width => 2,
      c_symmetry => 1,
      c_xdevicefamily => "artix7",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_15ffe94f3ff4129f
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tuser => s_axis_data_tuser,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tdata => m_axis_data_tdata,
    event_s_data_chanid_incorrect => event_s_data_chanid_incorrect
  );
-- synthesis translate_on

END fr_cmplr_v6_3_15ffe94f3ff4129f_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_2b018066c9a0cd8a.vhd when simulating
-- the core, fr_cmplr_v6_3_2b018066c9a0cd8a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_2b018066c9a0cd8a IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END fr_cmplr_v6_3_2b018066c9a0cd8a;

ARCHITECTURE fr_cmplr_v6_3_2b018066c9a0cd8a_a OF fr_cmplr_v6_3_2b018066c9a0cd8a IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_2b018066c9a0cd8a
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(47 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_2b018066c9a0cd8a USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "45,45",
      c_accum_path_widths => "45,45",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_2b018066c9a0cd8a.mif",
      c_coef_file_lines => 140,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0,0",
      c_coef_path_src => "0,0",
      c_coef_path_widths => "16,16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "4",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_2b018066c9a0cd8a",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 1,
      c_data_memtype => 1,
      c_data_path_sign => "0,0",
      c_data_path_src => "0,1",
      c_data_path_widths => "24,24",
      c_data_width => 24,
      c_datapath_memtype => 1,
      c_decim_rate => 35,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 12,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 1,
      c_m_data_tdata_width => 64,
      c_m_data_tuser_width => 1,
      c_mem_arrangement => 1,
      c_num_channels => 2,
      c_num_filts => 1,
      c_num_madds => 4,
      c_num_reload_slots => 1,
      c_num_taps => 248,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "25,25",
      c_output_rate => 35,
      c_output_width => 25,
      c_oversampling_rate => 1,
      c_reload_tdata_width => 1,
      c_round_mode => 4,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 1,
      c_s_data_tdata_width => 48,
      c_s_data_tuser_width => 1,
      c_symmetry => 1,
      c_xdevicefamily => "artix7",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_2b018066c9a0cd8a
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tuser => s_axis_data_tuser,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tdata => m_axis_data_tdata,
    event_s_data_chanid_incorrect => event_s_data_chanid_incorrect
  );
-- synthesis translate_on

END fr_cmplr_v6_3_2b018066c9a0cd8a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_8e79a078fc118dc6.vhd when simulating
-- the core, fr_cmplr_v6_3_8e79a078fc118dc6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_8e79a078fc118dc6 IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END fr_cmplr_v6_3_8e79a078fc118dc6;

ARCHITECTURE fr_cmplr_v6_3_8e79a078fc118dc6_a OF fr_cmplr_v6_3_8e79a078fc118dc6 IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_8e79a078fc118dc6
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_8e79a078fc118dc6 USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "42",
      c_accum_path_widths => "42",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_8e79a078fc118dc6.mif",
      c_coef_file_lines => 18,
      c_coef_mem_packing => 0,
      c_coef_memtype => 2,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "1",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_8e79a078fc118dc6",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 1,
      c_data_memtype => 1,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "24",
      c_data_width => 24,
      c_datapath_memtype => 2,
      c_decim_rate => 2,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 1400000,
      c_interp_rate => 1,
      c_ipbuff_memtype => 2,
      c_latency => 18,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 1,
      c_m_data_tdata_width => 32,
      c_m_data_tuser_width => 2,
      c_mem_arrangement => 1,
      c_num_channels => 4,
      c_num_filts => 1,
      c_num_madds => 1,
      c_num_reload_slots => 1,
      c_num_taps => 35,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "25",
      c_output_rate => 2800000,
      c_output_width => 25,
      c_oversampling_rate => 9,
      c_reload_tdata_width => 1,
      c_round_mode => 4,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 1,
      c_s_data_tdata_width => 24,
      c_s_data_tuser_width => 2,
      c_symmetry => 1,
      c_xdevicefamily => "artix7",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_8e79a078fc118dc6
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tuser => s_axis_data_tuser,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tdata => m_axis_data_tdata,
    event_s_data_chanid_incorrect => event_s_data_chanid_incorrect
  );
-- synthesis translate_on

END fr_cmplr_v6_3_8e79a078fc118dc6_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fr_cmplr_v6_3_b1697e0c92d2e32a.vhd when simulating
-- the core, fr_cmplr_v6_3_b1697e0c92d2e32a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fr_cmplr_v6_3_b1697e0c92d2e32a IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END fr_cmplr_v6_3_b1697e0c92d2e32a;

ARCHITECTURE fr_cmplr_v6_3_b1697e0c92d2e32a_a OF fr_cmplr_v6_3_b1697e0c92d2e32a IS
-- synthesis translate_off
COMPONENT wrapped_fr_cmplr_v6_3_b1697e0c92d2e32a
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tuser : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    event_s_data_chanid_incorrect : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fr_cmplr_v6_3_b1697e0c92d2e32a USE ENTITY XilinxCoreLib.fir_compiler_v6_3(behavioral)
    GENERIC MAP (
      c_accum_op_path_widths => "44",
      c_accum_path_widths => "44",
      c_channel_pattern => "fixed",
      c_coef_file => "fr_cmplr_v6_3_b1697e0c92d2e32a.mif",
      c_coef_file_lines => 240,
      c_coef_mem_packing => 0,
      c_coef_memtype => 1,
      c_coef_path_sign => "0",
      c_coef_path_src => "0",
      c_coef_path_widths => "16",
      c_coef_reload => 0,
      c_coef_width => 16,
      c_col_config => "1",
      c_col_mode => 1,
      c_col_pipe_len => 4,
      c_component_name => "fr_cmplr_v6_3_b1697e0c92d2e32a",
      c_config_packet_size => 0,
      c_config_sync_mode => 0,
      c_config_tdata_width => 1,
      c_data_has_tlast => 0,
      c_data_mem_packing => 0,
      c_data_memtype => 1,
      c_data_path_sign => "0",
      c_data_path_src => "0",
      c_data_path_widths => "25",
      c_data_width => 25,
      c_datapath_memtype => 2,
      c_decim_rate => 10,
      c_ext_mult_cnfg => "none",
      c_filter_type => 1,
      c_filts_packed => 0,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_config_channel => 0,
      c_input_rate => 5600000,
      c_interp_rate => 1,
      c_ipbuff_memtype => 0,
      c_latency => 31,
      c_m_data_has_tready => 0,
      c_m_data_has_tuser => 1,
      c_m_data_tdata_width => 32,
      c_m_data_tuser_width => 2,
      c_mem_arrangement => 0,
      c_num_channels => 4,
      c_num_filts => 1,
      c_num_madds => 1,
      c_num_reload_slots => 1,
      c_num_taps => 240,
      c_opbuff_memtype => 0,
      c_opt_madds => "none",
      c_optimization => 0,
      c_output_path_widths => "26",
      c_output_rate => 56000000,
      c_output_width => 26,
      c_oversampling_rate => 24,
      c_reload_tdata_width => 1,
      c_round_mode => 4,
      c_s_data_has_fifo => 0,
      c_s_data_has_tuser => 1,
      c_s_data_tdata_width => 32,
      c_s_data_tuser_width => 2,
      c_symmetry => 0,
      c_xdevicefamily => "artix7",
      c_zero_packing_factor => 1
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fr_cmplr_v6_3_b1697e0c92d2e32a
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tuser => s_axis_data_tuser,
    s_axis_data_tdata => s_axis_data_tdata,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tdata => m_axis_data_tdata,
    event_s_data_chanid_incorrect => event_s_data_chanid_incorrect
  );
-- synthesis translate_on

END fr_cmplr_v6_3_b1697e0c92d2e32a_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_7786f9df1b07f80e.vhd when simulating
-- the core, mult_11_2_7786f9df1b07f80e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_7786f9df1b07f80e IS
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(49 DOWNTO 0)
  );
END mult_11_2_7786f9df1b07f80e;

ARCHITECTURE mult_11_2_7786f9df1b07f80e_a OF mult_11_2_7786f9df1b07f80e IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_7786f9df1b07f80e
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(24 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(49 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_7786f9df1b07f80e USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_value => "10000001",
      c_b_width => 25,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 1,
      c_has_ce => 1,
      c_has_sclr => 1,
      c_has_zero_detect => 0,
      c_latency => 8,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 49,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "artix7"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_7786f9df1b07f80e
  PORT MAP (
    clk => clk,
    a => a,
    b => b,
    ce => ce,
    sclr => sclr,
    p => p
  );
-- synthesis translate_on

END mult_11_2_7786f9df1b07f80e_a;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlclockenablegenerator is
  generic (
    period: integer := 2;
    log_2_period: integer := 0;
    pipeline_regs: integer := 5
  );
  port (
    clk: in std_logic;
    clr: in std_logic;
    ce: out std_logic
  );
end xlclockenablegenerator;
architecture behavior of xlclockenablegenerator is
  component synth_reg_w_init
    generic (
      width: integer;
      init_index: integer;
      init_value: bit_vector;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function size_of_uint(inp: integer; power_of_2: boolean)
    return integer
  is
    constant inp_vec: std_logic_vector(31 downto 0) :=
      integer_to_std_logic_vector(inp,32, xlUnsigned);
    variable result: integer;
  begin
    result := 32;
    for i in 0 to 31 loop
      if inp_vec(i) = '1' then
        result := i;
      end if;
    end loop;
    if power_of_2 then
      return result;
    else
      return result+1;
    end if;
  end;
  function is_power_of_2(inp: std_logic_vector)
    return boolean
  is
    constant width: integer := inp'length;
    variable vec: std_logic_vector(width - 1 downto 0);
    variable single_bit_set: boolean;
    variable more_than_one_bit_set: boolean;
    variable result: boolean;
  begin
    vec := inp;
    single_bit_set := false;
    more_than_one_bit_set := false;
    -- synopsys translate_off
    if (is_XorU(vec)) then
      return false;
    end if;
     -- synopsys translate_on
    if width > 0 then
      for i in 0 to width - 1 loop
        if vec(i) = '1' then
          if single_bit_set then
            more_than_one_bit_set := true;
          end if;
          single_bit_set := true;
        end if;
      end loop;
    end if;
    if (single_bit_set and not(more_than_one_bit_set)) then
      result := true;
    else
      result := false;
    end if;
    return result;
  end;
  function ce_reg_init_val(index, period : integer)
    return integer
  is
     variable result: integer;
   begin
      result := 0;
      if ((index mod period) = 0) then
          result := 1;
      end if;
      return result;
  end;
  function remaining_pipe_regs(num_pipeline_regs, period : integer)
    return integer
  is
     variable factor, result: integer;
  begin
      factor := (num_pipeline_regs / period);
      result := num_pipeline_regs - (period * factor) + 1;
      return result;
  end;

  function sg_min(L, R: INTEGER) return INTEGER is
  begin
      if L < R then
            return L;
      else
            return R;
      end if;
  end;
  constant max_pipeline_regs : integer := 8;
  constant pipe_regs : integer := 5;
  constant num_pipeline_regs : integer := sg_min(pipeline_regs, max_pipeline_regs);
  constant rem_pipeline_regs : integer := remaining_pipe_regs(num_pipeline_regs,period);
  constant period_floor: integer := max(2, period);
  constant power_of_2_counter: boolean :=
    is_power_of_2(integer_to_std_logic_vector(period_floor,32, xlUnsigned));
  constant cnt_width: integer :=
    size_of_uint(period_floor, power_of_2_counter);
  constant clk_for_ce_pulse_minus1: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector((period_floor - 2),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus2: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - 3),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus_regs: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - rem_pipeline_regs),cnt_width, xlUnsigned);
  signal clk_num: unsigned(cnt_width - 1 downto 0) := (others => '0');
  signal ce_vec : std_logic_vector(num_pipeline_regs downto 0);
  signal internal_ce: std_logic_vector(0 downto 0);
  signal cnt_clr, cnt_clr_dly: std_logic_vector (0 downto 0);
begin
  cntr_gen: process(clk)
  begin
    if clk'event and clk = '1'  then
        if ((cnt_clr_dly(0) = '1') or (clr = '1')) then
          clk_num <= (others => '0');
        else
          clk_num <= clk_num + 1;
        end if;
    end if;
  end process;
  clr_gen: process(clk_num, clr)
  begin
    if power_of_2_counter then
      cnt_clr(0) <= clr;
    else
      if (unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus1
          or clr = '1') then
        cnt_clr(0) <= '1';
      else
        cnt_clr(0) <= '0';
      end if;
    end if;
  end process;
  clr_reg: synth_reg_w_init
    generic map (
      width => 1,
      init_index => 0,
      init_value => b"0000",
      latency => 1
    )
    port map (
      i => cnt_clr,
      ce => '1',
      clr => clr,
      clk => clk,
      o => cnt_clr_dly
    );
  pipelined_ce : if period > 1 generate
      ce_gen: process(clk_num)
      begin
          if unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus_regs then
              ce_vec(num_pipeline_regs) <= '1';
          else
              ce_vec(num_pipeline_regs) <= '0';
          end if;
      end process;
      ce_pipeline: for index in num_pipeline_regs downto 1 generate
          ce_reg : synth_reg_w_init
              generic map (
                  width => 1,
                  init_index => ce_reg_init_val(index, period),
                  init_value => b"0000",
                  latency => 1
                  )
              port map (
                  i => ce_vec(index downto index),
                  ce => '1',
                  clr => clr,
                  clk => clk,
                  o => ce_vec(index-1 downto index-1)
                  );
      end generate;
      internal_ce <= ce_vec(0 downto 0);
  end generate;
  generate_clock_enable: if period > 1 generate
    ce <= internal_ce(0);
  end generate;
  generate_clock_enable_constant: if period = 1 generate
    ce <= '1';
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_cd3162dc0d is
  port (
    in0 : in std_logic_vector((16 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_cd3162dc0d;


architecture behavior of concat_cd3162dc0d is
  signal in0_1_23: unsigned((16 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((24 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_91ef1678ca is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_91ef1678ca;


architecture behavior of constant_91ef1678ca is
begin
  op <= "00000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_7025463ea8 is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_7025463ea8;


architecture behavior of reinterpret_7025463ea8 is
  signal input_port_1_40: signed((16 - 1) downto 0);
  signal output_port_5_5_force: unsigned((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_f21e7f2ddf is
  port (
    input_port : in std_logic_vector((8 - 1) downto 0);
    output_port : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_f21e7f2ddf;


architecture behavior of reinterpret_f21e7f2ddf is
  signal input_port_1_40: unsigned((8 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_4bf1ad328a is
  port (
    input_port : in std_logic_vector((24 - 1) downto 0);
    output_port : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_4bf1ad328a;


architecture behavior of reinterpret_4bf1ad328a is
  signal input_port_1_40: unsigned((24 - 1) downto 0);
  signal output_port_5_5_force: signed((24 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlceprobe is
    generic (d_width  : integer := 8;
             q_width  : integer := 1);
    port (d       : in std_logic_vector (d_width-1 downto 0);
          ce      : in std_logic;
          clk     : in std_logic;
          q       : out std_logic_vector (q_width-1 downto 0));
end xlceprobe;
architecture behavior of xlceprobe is
    component BUF
        port(
            O  :        out   STD_ULOGIC;
            I  :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of BUF : component is true;
    attribute fpga_dont_touch of BUF : component is "true";
    signal ce_vec : std_logic_vector(0 downto 0);
begin
    buf_comp : buf port map(i => ce, o => ce_vec(0));
    q <= ce_vec;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_a2121d82da is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((24 - 1) downto 0);
    d1 : in std_logic_vector((24 - 1) downto 0);
    y : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_a2121d82da;


architecture behavior of mux_a2121d82da is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((24 - 1) downto 0);
  signal d1_1_27: std_logic_vector((24 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((24 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity counter_41314d726b is
  port (
    rst : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end counter_41314d726b;


architecture behavior of counter_41314d726b is
  signal rst_1_40: boolean;
  signal en_1_45: boolean;
  signal count_reg_20_23: unsigned((1 - 1) downto 0) := "0";
  signal count_reg_20_23_rst: std_logic;
  signal count_reg_20_23_en: std_logic;
  signal bool_44_4: boolean;
  signal rst_limit_join_44_1: boolean;
  signal count_reg_join_44_1: unsigned((2 - 1) downto 0);
  signal count_reg_join_44_1_en: std_logic;
  signal count_reg_join_44_1_rst: std_logic;
begin
  rst_1_40 <= ((rst) = "1");
  en_1_45 <= ((en) = "1");
  proc_count_reg_20_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (count_reg_20_23_rst = '1')) then
        count_reg_20_23 <= "0";
      elsif ((ce = '1') and (count_reg_20_23_en = '1')) then
        count_reg_20_23 <= count_reg_20_23 + std_logic_vector_to_unsigned("1");
      end if;
    end if;
  end process proc_count_reg_20_23;
  bool_44_4 <= rst_1_40 or false;
  proc_if_44_1: process (bool_44_4, count_reg_20_23, en_1_45)
  is
  begin
    if bool_44_4 then
      count_reg_join_44_1_rst <= '1';
    elsif en_1_45 then
      count_reg_join_44_1_rst <= '0';
    else
      count_reg_join_44_1_rst <= '0';
    end if;
    if en_1_45 then
      count_reg_join_44_1_en <= '1';
    else
      count_reg_join_44_1_en <= '0';
    end if;
    if bool_44_4 then
      rst_limit_join_44_1 <= false;
    elsif en_1_45 then
      rst_limit_join_44_1 <= false;
    else
      rst_limit_join_44_1 <= false;
    end if;
  end process proc_if_44_1;
  count_reg_20_23_rst <= count_reg_join_44_1_rst;
  count_reg_20_23_en <= count_reg_join_44_1_en;
  op <= unsigned_to_std_logic_vector(count_reg_20_23);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlusamp is
    generic (
             d_width      : integer := 5;
             d_bin_pt     : integer := 2;
             d_arith      : integer := xlUnsigned;
             q_width      : integer := 5;
             q_bin_pt     : integer := 2;
             q_arith      : integer := xlUnsigned;
             en_width     : integer := 1;
             en_bin_pt    : integer := 0;
             en_arith     : integer := xlUnsigned;
             sampling_ratio     : integer := 2;
             latency      : integer := 1;
             copy_samples : integer := 0);
    port (
          d        : in std_logic_vector (d_width-1 downto 0);
          src_clk  : in std_logic;
          src_ce   : in std_logic;
          src_clr  : in std_logic;
          dest_clk : in std_logic;
          dest_ce  : in std_logic;
          dest_clr : in std_logic;
          en       : in std_logic_vector(en_width-1 downto 0);
          q        : out std_logic_vector (q_width-1 downto 0)
         );
end xlusamp;
architecture struct of xlusamp is
    component synth_reg
      generic (
        width: integer := 16;
        latency: integer := 5
      );
      port (
        i: in std_logic_vector(width - 1 downto 0);
        ce: in std_logic;
        clr: in std_logic;
        clk: in std_logic;
        o: out std_logic_vector(width - 1 downto 0)
      );
    end component;
    component FDSE
        port (q  : out   std_ulogic;
              d  : in    std_ulogic;
              c  : in    std_ulogic;
              s  : in    std_ulogic;
              ce : in    std_ulogic);
    end component;
    attribute syn_black_box of FDSE : component is true;
    attribute fpga_dont_touch of FDSE : component is "true";
    signal zero    : std_logic_vector (d_width-1 downto 0);
    signal mux_sel : std_logic;
    signal sampled_d  : std_logic_vector (d_width-1 downto 0);
    signal internal_ce : std_logic;
begin
   sel_gen : FDSE
                port map (q  => mux_sel,
                        d  => src_ce,
            c  => src_clk,
            s  => src_clr,
            ce => dest_ce);
  internal_ce <= src_ce and en(0);
  copy_samples_false : if (copy_samples = 0) generate
      zero <= (others => '0');
      gen_q_cp_smpls_0_and_lat_0: if (latency = 0) generate
        cp_smpls_0_and_lat_0: process (mux_sel, d, zero)
        begin
          if (mux_sel = '1') then
            q <= d;
          else
            q <= zero;
          end if;
        end process cp_smpls_0_and_lat_0;
      end generate;
      gen_q_cp_smpls_0_and_lat_gt_0: if (latency > 0) generate
        sampled_d_reg: synth_reg
          generic map (
            width => d_width,
            latency => latency
          )
          port map (
            i => d,
            ce => internal_ce,
            clr => src_clr,
            clk => src_clk,
            o => sampled_d
          );

        gen_q_check_mux_sel: process (mux_sel, sampled_d, zero)
        begin
          if (mux_sel = '1') then
            q <= sampled_d;
          else
            q <= zero;
          end if;
        end process gen_q_check_mux_sel;
      end generate;
   end generate;
   copy_samples_true : if (copy_samples = 1) generate
     gen_q_cp_smpls_1_and_lat_0: if (latency = 0) generate
       q <= d;
     end generate;
     gen_q_cp_smpls_1_and_lat_gt_0: if (latency > 0) generate
       q <= sampled_d;
       sampled_d_reg2: synth_reg
         generic map (
           width => d_width,
           latency => latency
         )
         port map (
           i => d,
           ce => internal_ce,
           clr => src_clr,
           clk => src_clk,
           o => sampled_d
         );
     end generate;
   end generate;
end architecture struct;
-------------------------------------------------------------------------------
-- Title      : Look-up table sweeper
-- Project    :
-------------------------------------------------------------------------------
-- File       : lut_sweep.vhd
-- Author     : aylons  <aylons@LNLS190>
-- Company    :
-- Created    : 2014-03-07
-- Last update: 2014-03-07
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Tool for sweeping through look-up table addresses
-------------------------------------------------------------------------------
-- Copyright (c) 2014
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-03-07  1.0      aylons  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

-------------------------------------------------------------------------------

entity lut_sweep is
  generic (
    g_bus_size      : natural := 8;
    g_first_address : natural := 0;
    g_last_address  : natural := 147;
    g_sweep_mode    : string  := "sawtooth"
    );
  port (
    rst_n_i   : in  std_logic;
    clk_i     : in  std_logic;
    ce_i      : in  std_logic;
    address_o : out std_logic_vector(g_bus_size-1 downto 0));
end entity lut_sweep;

-------------------------------------------------------------------------------

architecture str of lut_sweep is

begin  -- architecture str

  counting : process(clk_i)
    variable count : natural := 0;
  begin

    if rising_edge(clk_i) then

      if rst_n_i = '0' then
        count        := 0;

      elsif ce_i = '1' then
        if count = g_last_address then
          count := g_first_address;
        else
          count := count + 1;
        end if;  --count = last_address

        address_o <= std_logic_vector(to_unsigned(count, g_bus_size));
      end if;  -- reset
    end if;  -- rising_edge

  end process counting;


end architecture str;

-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Title      : Fixed sin-cos DDS
-- Project    :
-------------------------------------------------------------------------------
-- File       : fixed_dds.vhd
-- Author     : aylons  <aylons@LNLS190>
-- Company    :
-- Created    : 2014-03-07
-- Last update: 2014-03-07
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Fixed frequency phase and quadrature DDS for use in tuned DDCs.
-------------------------------------------------------------------------------
-- Copyright (c) 2014
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2014-03-07  1.0      aylons  Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

library work;
use work.genram_pkg.all;
-------------------------------------------------------------------------------

entity fixed_dds is

  generic (
    g_number_of_points : natural := 148;
    g_output_width     : natural := 24;
    g_dither           : boolean := false;
    g_sin_file         : string  := "./dds_sin.ram";
    g_cos_file         : string  := "./dds_cos.ram"
    );
  port (
    clk_i     : in  std_logic;
    ce_i      : in  std_logic;
    rst_n_i   : in  std_logic;
    sin_o     : out std_logic_vector(g_output_width-1 downto 0);
    cos_o     : out std_logic_vector(g_output_width-1 downto 0)
    );

end entity fixed_dds;

-------------------------------------------------------------------------------

architecture str of fixed_dds is

  constant c_bus_size : natural := f_log2_size(g_number_of_points);
  signal cur_address  : std_logic_vector(c_bus_size-1 downto 0);

  component generic_simple_dpram is
    generic (
      g_data_width               : natural;
      g_size                     : natural;
      g_with_byte_enable         : boolean;
      g_addr_conflict_resolution : string;
      g_init_file                : string;
      g_dual_clock               : boolean);
    port (
      rst_n_i : in  std_logic                                        := '1';
      clka_i  : in  std_logic;
      bwea_i  : in  std_logic_vector((g_data_width+7)/8 -1 downto 0) := f_gen_dummy_vec('1', (g_data_width+7)/8);
      wea_i   : in  std_logic;
      aa_i    : in  std_logic_vector(c_bus_size-1 downto 0);
      da_i    : in  std_logic_vector(g_data_width-1 downto 0);
      clkb_i  : in  std_logic;
      ab_i    : in  std_logic_vector(c_bus_size-1 downto 0);
      qb_o    : out std_logic_vector(g_data_width-1 downto 0));
  end component generic_simple_dpram;

  component lut_sweep is
    generic (
      g_bus_size      : natural;
      g_first_address : natural;
      g_last_address  : natural;
      g_sweep_mode    : string);
    port (
      rst_n_i : in  std_logic;
      clk_i   : in  std_logic;
      ce_i      : in  std_logic;
      address_o : out std_logic_vector(c_bus_size-1 downto 0));
  end component lut_sweep;

begin  -- architecture str

  cmp_sin_lut : generic_simple_dpram
    generic map (
      g_data_width               => g_output_width,
      g_size                     => g_number_of_points,
      g_with_byte_enable         => false,
      g_addr_conflict_resolution => "dont_care",
      g_init_file                => g_sin_file,
      g_dual_clock               => false
      )
    port map (
      rst_n_i => rst_n_i,
      clka_i  => clk_i,
      bwea_i  => (others => '0'),
      wea_i   => '0',
      aa_i    => cur_address,
      da_i    => (others => '0'),
      clkb_i  => clk_i,
      ab_i    => cur_address,
      qb_o    => sin_o
      );

  cmp_cos_lut : generic_simple_dpram
    generic map (
      g_data_width               => g_output_width,
      g_size                     => g_number_of_points,
      g_with_byte_enable         => false,
      g_addr_conflict_resolution => "dont_care",
      g_init_file                => g_cos_file,
      g_dual_clock               => false
      )
    port map (
      rst_n_i => rst_n_i,
      clka_i  => clk_i,
      bwea_i  => (others => '0'),
      wea_i   => '0',
      aa_i    => cur_address,
      da_i    => (others => '0'),
      clkb_i  => clk_i,
      ab_i    => cur_address,
      qb_o    => cos_o
      );

  cmp_sweep : lut_sweep
    generic map (
      g_bus_size      => c_bus_size,
      g_first_address => 0,
      g_last_address  => g_number_of_points-1,
      g_sweep_mode    => "sawtooth")
    port map (
      rst_n_i => rst_n_i,
      clk_i   => clk_i,
      ce_i      => ce_i,
      address_o => cur_address);

end architecture str;

-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xldsamp is
  generic (
    d_width: integer := 12;
    d_bin_pt: integer := 0;
    d_arith: integer := xlUnsigned;
    q_width: integer := 12;
    q_bin_pt: integer := 0;
    q_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    ds_ratio: integer := 2;
    phase: integer := 0;
    latency: integer := 1
  );
  port (
    d: in std_logic_vector(d_width - 1 downto 0);
    src_clk: in std_logic;
    src_ce: in std_logic;
    src_clr: in std_logic;
    dest_clk: in std_logic;
    dest_ce: in std_logic;
    dest_clr: in std_logic;
    en: in std_logic_vector(en_width - 1 downto 0);
    q: out std_logic_vector(q_width - 1 downto 0)
  );
end xldsamp;
architecture struct of xldsamp is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component fdse
    port (
      q: out   std_ulogic;
      d: in    std_ulogic;
      c: in    std_ulogic;
      s: in    std_ulogic;
      ce: in    std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  signal adjusted_dest_ce: std_logic;
  signal adjusted_dest_ce_w_en: std_logic;
  signal dest_ce_w_en: std_logic;
  signal smpld_d: std_logic_vector(d_width-1 downto 0);
begin
  adjusted_ce_needed: if ((latency = 0) or (phase /= (ds_ratio - 1))) generate
    dest_ce_reg: fdse
      port map (
        q => adjusted_dest_ce,
        d => dest_ce,
        c => src_clk,
        s => src_clr,
        ce => src_ce
      );
  end generate;
  latency_eq_0: if (latency = 0) generate
    shutter_d_reg: synth_reg
      generic map (
        width => d_width,
        latency => 1
      )
      port map (
        i => d,
        ce => adjusted_dest_ce,
        clr => src_clr,
        clk => src_clk,
        o => smpld_d
      );
    shutter_mux: process (adjusted_dest_ce, d, smpld_d)
    begin
      if adjusted_dest_ce = '0' then
        q <= smpld_d;
      else
        q <= d;
      end if;
    end process;
  end generate;
  latency_gt_0: if (latency > 0) generate
    dbl_reg_test: if (phase /= (ds_ratio-1)) generate
        smpl_d_reg: synth_reg
          generic map (
            width => d_width,
            latency => 1
          )
          port map (
            i => d,
            ce => adjusted_dest_ce_w_en,
            clr => src_clr,
            clk => src_clk,
            o => smpld_d
          );
    end generate;
    sngl_reg_test: if (phase = (ds_ratio -1)) generate
      smpld_d <= d;
    end generate;
    latency_pipe: synth_reg
      generic map (
        width => d_width,
        latency => latency
      )
      port map (
        i => smpld_d,
        ce => dest_ce_w_en,
        clr => src_clr,
        clk => dest_clk,
        o => q
      );
  end generate;
  dest_ce_w_en <= dest_ce and en(0);
  adjusted_dest_ce_w_en <= adjusted_dest_ce and en(0);
end architecture struct;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_a892e1bf40 is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_a892e1bf40;


architecture behavior of relational_a892e1bf40 is
  signal a_1_31: unsigned((1 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  type array_type_op_mem_32_22 is array (0 to (1 - 1)) of boolean;
  signal op_mem_32_22: array_type_op_mem_32_22 := (
    0 => false);
  signal op_mem_32_22_front_din: boolean;
  signal op_mem_32_22_back: boolean;
  signal op_mem_32_22_push_front_pop_back_en: std_logic;
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  op_mem_32_22_back <= op_mem_32_22(0);
  proc_op_mem_32_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_32_22_push_front_pop_back_en = '1')) then
        op_mem_32_22(0) <= op_mem_32_22_front_din;
      end if;
    end if;
  end process proc_op_mem_32_22;
  result_12_3_rel <= a_1_31 = b_1_34;
  op_mem_32_22_front_din <= result_12_3_rel;
  op_mem_32_22_push_front_pop_back_en <= '1';
  op <= boolean_to_vector(op_mem_32_22_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_b62f4240f0 is
  port (
    input_port : in std_logic_vector((24 - 1) downto 0);
    output_port : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_b62f4240f0;


architecture behavior of reinterpret_b62f4240f0 is
  signal input_port_1_40: signed((24 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcordic_3fb964e2f71602f328fdd11ab57d7304 is
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_phase:out std_logic_vector(23 downto 0);
    m_axis_dout_tdata_real:out std_logic_vector(23 downto 0);
    m_axis_dout_tuser_cartesian_tuser:out std_logic_vector(0 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_cartesian_tdata_imag:in std_logic_vector(24 downto 0);
    s_axis_cartesian_tdata_real:in std_logic_vector(24 downto 0);
    s_axis_cartesian_tuser_user:in std_logic_vector(0 downto 0);
    s_axis_cartesian_tvalid:in std_logic
  );
end xlcordic_3fb964e2f71602f328fdd11ab57d7304;


architecture behavior of xlcordic_3fb964e2f71602f328fdd11ab57d7304  is
  component crdc_v5_0_3d2446e74ce31176
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(47 downto 0);
      m_axis_dout_tuser:out std_logic_vector(0 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_cartesian_tdata:in std_logic_vector(63 downto 0);
      s_axis_cartesian_tuser:in std_logic_vector(0 downto 0);
      s_axis_cartesian_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal m_axis_dout_tuser_net: std_logic_vector(0 downto 0) := (others=>'0');
signal s_axis_cartesian_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
signal s_axis_cartesian_tuser_net: std_logic_vector(0 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_phase <= m_axis_dout_tdata_net(47 downto 24);
  m_axis_dout_tdata_real <= m_axis_dout_tdata_net(23 downto 0);
  m_axis_dout_tuser_cartesian_tuser <= m_axis_dout_tuser_net(0 downto 0);
  s_axis_cartesian_tdata_net(56 downto 32) <= s_axis_cartesian_tdata_imag;
  s_axis_cartesian_tdata_net(24 downto 0) <= s_axis_cartesian_tdata_real;
  s_axis_cartesian_tuser_net(0 downto 0) <= s_axis_cartesian_tuser_user;
  crdc_v5_0_3d2446e74ce31176_instance : crdc_v5_0_3d2446e74ce31176
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tuser=>m_axis_dout_tuser_net,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_cartesian_tdata=>s_axis_cartesian_tdata_net,
      s_axis_cartesian_tuser=>s_axis_cartesian_tuser_net,
      s_axis_cartesian_tvalid=>s_axis_cartesian_tvalid
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_31a4235b32 is
  port (
    input_port : in std_logic_vector((25 - 1) downto 0);
    output_port : out std_logic_vector((25 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_31a4235b32;


architecture behavior of reinterpret_31a4235b32 is
  signal input_port_1_40: signed((25 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_fa01b5fd95 is
  port (
    input_port : in std_logic_vector((58 - 1) downto 0);
    output_port : out std_logic_vector((58 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_fa01b5fd95;


architecture behavior of reinterpret_fa01b5fd95 is
  signal input_port_1_40: signed((58 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cda50df78a is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cda50df78a;


architecture behavior of constant_cda50df78a is
begin
  op <= "00";
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer :=  0;
           reset        : integer :=  0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        rst     : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if ((reg_retiming = 0) and (reset = 0)) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if ((reg_retiming = 1) or (reset = 1)) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => rst,
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_d29d27b7b3 is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_d29d27b7b3;


architecture behavior of relational_d29d27b7b3 is
  signal a_1_31: unsigned((1 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  type array_type_op_mem_32_22 is array (0 to (1 - 1)) of boolean;
  signal op_mem_32_22: array_type_op_mem_32_22 := (
    0 => false);
  signal op_mem_32_22_front_din: boolean;
  signal op_mem_32_22_back: boolean;
  signal op_mem_32_22_push_front_pop_back_en: std_logic;
  signal cast_12_12: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  op_mem_32_22_back <= op_mem_32_22(0);
  proc_op_mem_32_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_32_22_push_front_pop_back_en = '1')) then
        op_mem_32_22(0) <= op_mem_32_22_front_din;
      end if;
    end if;
  end process proc_op_mem_32_22;
  cast_12_12 <= u2u_cast(a_1_31, 0, 2, 0);
  result_12_3_rel <= cast_12_12 = b_1_34;
  op_mem_32_22_front_din <= result_12_3_rel;
  op_mem_32_22_push_front_pop_back_en <= '1';
  op <= boolean_to_vector(op_mem_32_22_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcic_compiler_2d3b496704eca3daaae85383d488a908 is
  port(
    ce:in std_logic;
    ce_1120:in std_logic;
    ce_logic_1:in std_logic;
    clk:in std_logic;
    clk_1120:in std_logic;
    clk_logic_1:in std_logic;
    event_tlast_missing:out std_logic;
    event_tlast_unexpected:out std_logic;
    m_axis_data_tdata_data:out std_logic_vector(57 downto 0);
    m_axis_data_tlast:out std_logic;
    m_axis_data_tuser_chan_out:out std_logic_vector(0 downto 0);
    m_axis_data_tuser_chan_sync:out std_logic_vector(0 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_data:in std_logic_vector(23 downto 0);
    s_axis_data_tlast:in std_logic;
    s_axis_data_tready:out std_logic
  );
end xlcic_compiler_2d3b496704eca3daaae85383d488a908;


architecture behavior of xlcic_compiler_2d3b496704eca3daaae85383d488a908  is
  component cc_cmplr_v3_0_964aa42461b15ac2
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_tlast_missing:out std_logic;
      event_tlast_unexpected:out std_logic;
      m_axis_data_tdata:out std_logic_vector(63 downto 0);
      m_axis_data_tlast:out std_logic;
      m_axis_data_tuser:out std_logic_vector(15 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tlast:in std_logic;
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net: std_logic_vector(57 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_captured: std_logic_vector(57 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_or_captured_net: std_logic_vector(57 downto 0) := (others=>'0');
signal m_axis_data_tlast_ps_net: std_logic := '0';
signal m_axis_data_tlast_ps_net_captured: std_logic := '0';
signal m_axis_data_tlast_ps_net_or_captured_net: std_logic := '0';
signal m_axis_data_tuser_net: std_logic_vector(15 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net_captured: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net_or_captured_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net_captured: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net_or_captured_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_data_ps_net <= m_axis_data_tdata_net(57 downto 0);
  m_axis_data_tuser_chan_sync_ps_net <= m_axis_data_tuser_net(8 downto 8);
  m_axis_data_tuser_chan_out_ps_net <= m_axis_data_tuser_net(0 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_data;
  m_axis_data_tdata_data_ps_net_or_captured_net <= m_axis_data_tdata_data_ps_net or m_axis_data_tdata_data_ps_net_captured;
m_axis_data_tdata_data_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 58,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net_or_captured_net,
        ce => ce_1120,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tdata_data
    );
m_axis_data_tdata_data_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 58,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tdata_data_ps_net_captured
    );
  m_axis_data_tlast_ps_net_or_captured_net <= m_axis_data_tlast_ps_net or m_axis_data_tlast_ps_net_captured;
m_axis_data_tlast_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tlast_ps_net_or_captured_net,
        ce => ce_1120,
        clr => '0',
        clk => clk_1120,
        o(0) => m_axis_data_tlast
    );
m_axis_data_tlast_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tlast_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1120,
        o(0) => m_axis_data_tlast_ps_net_captured
    );
  m_axis_data_tuser_chan_sync_ps_net_or_captured_net <= m_axis_data_tuser_chan_sync_ps_net or m_axis_data_tuser_chan_sync_ps_net_captured;
m_axis_data_tuser_chan_sync_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_sync_ps_net_or_captured_net,
        ce => ce_1120,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tuser_chan_sync
    );
m_axis_data_tuser_chan_sync_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_sync_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tuser_chan_sync_ps_net_captured
    );
  m_axis_data_tuser_chan_out_ps_net_or_captured_net <= m_axis_data_tuser_chan_out_ps_net or m_axis_data_tuser_chan_out_ps_net_captured;
m_axis_data_tuser_chan_out_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_out_ps_net_or_captured_net,
        ce => ce_1120,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tuser_chan_out
    );
m_axis_data_tuser_chan_out_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_out_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1120,
        o => m_axis_data_tuser_chan_out_ps_net_captured
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_1120,
        clr => '0',
        clk => clk_1120,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1120,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  cc_cmplr_v3_0_964aa42461b15ac2_instance : cc_cmplr_v3_0_964aa42461b15ac2
    port map(
      aclk=>clk,
      aclken=>ce,
      event_tlast_missing=>event_tlast_missing,
      event_tlast_unexpected=>event_tlast_unexpected,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tlast=>m_axis_data_tlast_ps_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tlast=>s_axis_data_tlast,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_1
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_9934b94a22 is
  port (
    input_port : in std_logic_vector((26 - 1) downto 0);
    output_port : out std_logic_vector((26 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_9934b94a22;


architecture behavior of reinterpret_9934b94a22 is
  signal input_port_1_40: unsigned((26 - 1) downto 0);
  signal output_port_5_5_force: signed((26 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlslice is
    generic (
        new_msb      : integer := 9;
        new_lsb      : integer := 1;
        x_width      : integer := 16;
        y_width      : integer := 8);
    port (
        x : in std_logic_vector (x_width-1 downto 0);
        y : out std_logic_vector (y_width-1 downto 0));
end xlslice;
architecture behavior of xlslice is
begin
    y <= x(new_msb downto new_lsb);
end  behavior;

-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlmult is
  generic (
    core_name0: string := "";
    a_width: integer := 4;
    a_bin_pt: integer := 2;
    a_arith: integer := xlSigned;
    b_width: integer := 4;
    b_bin_pt: integer := 1;
    b_arith: integer := xlSigned;
    p_width: integer := 8;
    p_bin_pt: integer := 2;
    p_arith: integer := xlSigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    extra_registers: integer := 0;
    c_a_width: integer := 7;
    c_b_width: integer := 7;
    c_type: integer := 0;
    c_a_type: integer := 0;
    c_b_type: integer := 0;
    c_pipelined: integer := 1;
    c_baat: integer := 4;
    multsign: integer := xlSigned;
    c_output_width: integer := 16
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    core_ce: in std_logic := '0';
    core_clr: in std_logic := '0';
    core_clk: in std_logic := '0';
    rst: in std_logic_vector(rst_width - 1 downto 0);
    en: in std_logic_vector(en_width - 1 downto 0);
    p: out std_logic_vector(p_width - 1 downto 0)
  );
end xlmult;
architecture behavior of xlmult is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component mult_11_2_7786f9df1b07f80e
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      clk: in std_logic;
      ce: in std_logic;
      sclr: in std_logic;
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of mult_11_2_7786f9df1b07f80e:
    component is true;
  attribute fpga_dont_touch of mult_11_2_7786f9df1b07f80e:
    component is "true";
  attribute box_type of mult_11_2_7786f9df1b07f80e:
    component  is "black_box";
  signal tmp_a: std_logic_vector(c_a_width - 1 downto 0);
  signal conv_a: std_logic_vector(c_a_width - 1 downto 0);
  signal tmp_b: std_logic_vector(c_b_width - 1 downto 0);
  signal conv_b: std_logic_vector(c_b_width - 1 downto 0);
  signal tmp_p: std_logic_vector(c_output_width - 1 downto 0);
  signal conv_p: std_logic_vector(p_width - 1 downto 0);
  -- synopsys translate_off
  signal real_a, real_b, real_p: real;
  -- synopsys translate_on
  signal rfd: std_logic;
  signal rdy: std_logic;
  signal nd: std_logic;
  signal internal_ce: std_logic;
  signal internal_clr: std_logic;
  signal internal_core_ce: std_logic;
begin
-- synopsys translate_off
-- synopsys translate_on
  internal_ce <= ce and en(0);
  internal_core_ce <= core_ce and en(0);
  internal_clr <= (clr or rst(0)) and ce;
  nd <= internal_ce;
  input_process:  process (a,b)
  begin
    tmp_a <= zero_ext(a, c_a_width);
    tmp_b <= zero_ext(b, c_b_width);
  end process;
  output_process: process (tmp_p)
  begin
    conv_p <= convert_type(tmp_p, c_output_width, a_bin_pt+b_bin_pt, multsign,
                           p_width, p_bin_pt, p_arith, quantization, overflow);
  end process;
  comp0: if ((core_name0 = "mult_11_2_7786f9df1b07f80e")) generate
    core_instance0: mult_11_2_7786f9df1b07f80e
      port map (
        a => tmp_a,
        clk => clk,
        ce => internal_ce,
        sclr => internal_clr,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  latency_gt_0: if (extra_registers > 0) generate
    reg: synth_reg
      generic map (
        width => p_width,
        latency => extra_registers
      )
      port map (
        i => conv_p,
        ce => internal_ce,
        clr => internal_clr,
        clk => clk,
        o => p
      );
  end generate;
  latency_eq_0: if (extra_registers = 0) generate
    p <= conv_p;
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcomplex_multiplier_456da30af0f77a480cf80f52b29b4396 is
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_imag:out std_logic_vector(23 downto 0);
    m_axis_dout_tdata_real:out std_logic_vector(23 downto 0);
    m_axis_dout_tuser:out std_logic_vector(0 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_a_tdata_imag:in std_logic_vector(23 downto 0);
    s_axis_a_tdata_real:in std_logic_vector(23 downto 0);
    s_axis_a_tvalid:in std_logic;
    s_axis_b_tdata_imag:in std_logic_vector(23 downto 0);
    s_axis_b_tdata_real:in std_logic_vector(23 downto 0);
    s_axis_b_tuser:in std_logic_vector(0 downto 0);
    s_axis_b_tvalid:in std_logic
  );
end xlcomplex_multiplier_456da30af0f77a480cf80f52b29b4396;


architecture behavior of xlcomplex_multiplier_456da30af0f77a480cf80f52b29b4396  is
  component cmpy_v5_0_02d02e0a23eb9773
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(47 downto 0);
      m_axis_dout_tuser:out std_logic_vector(0 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_a_tdata:in std_logic_vector(47 downto 0);
      s_axis_a_tvalid:in std_logic;
      s_axis_b_tdata:in std_logic_vector(47 downto 0);
      s_axis_b_tuser:in std_logic_vector(0 downto 0);
      s_axis_b_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal s_axis_a_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal s_axis_b_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_imag <= m_axis_dout_tdata_net(47 downto 24);
  m_axis_dout_tdata_real <= m_axis_dout_tdata_net(23 downto 0);
  s_axis_a_tdata_net(47 downto 24) <= s_axis_a_tdata_imag;
  s_axis_a_tdata_net(23 downto 0) <= s_axis_a_tdata_real;
  s_axis_b_tdata_net(47 downto 24) <= s_axis_b_tdata_imag;
  s_axis_b_tdata_net(23 downto 0) <= s_axis_b_tdata_real;
  cmpy_v5_0_02d02e0a23eb9773_instance : cmpy_v5_0_02d02e0a23eb9773
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tuser=>m_axis_dout_tuser,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_a_tdata=>s_axis_a_tdata_net,
      s_axis_a_tvalid=>s_axis_a_tvalid,
      s_axis_b_tdata=>s_axis_b_tdata_net,
      s_axis_b_tuser=>s_axis_b_tuser,
      s_axis_b_tvalid=>s_axis_b_tvalid
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_961b43f67a is
  port (
    d : in std_logic_vector((24 - 1) downto 0);
    q : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_961b43f67a;


architecture behavior of delay_961b43f67a is
  signal d_1_22: std_logic_vector((24 - 1) downto 0);
begin
  d_1_22 <= d;
  q <= d_1_22;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_f394f3309c is
  port (
    op : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_f394f3309c;


architecture behavior of constant_f394f3309c is
begin
  op <= "000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_c88e29aa6b is
  port (
    input_port : in std_logic_vector((61 - 1) downto 0);
    output_port : out std_logic_vector((61 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_c88e29aa6b;


architecture behavior of reinterpret_c88e29aa6b is
  signal input_port_1_40: signed((61 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_3a9a3daeb9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_3a9a3daeb9;


architecture behavior of constant_3a9a3daeb9 is
begin
  op <= "11";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a7e2bb9e12 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a7e2bb9e12;


architecture behavior of constant_a7e2bb9e12 is
begin
  op <= "01";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e8ddc079e9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e8ddc079e9;


architecture behavior of constant_e8ddc079e9 is
begin
  op <= "10";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_367321bc0c is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_367321bc0c;


architecture behavior of relational_367321bc0c is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  type array_type_op_mem_32_22 is array (0 to (1 - 1)) of boolean;
  signal op_mem_32_22: array_type_op_mem_32_22 := (
    0 => false);
  signal op_mem_32_22_front_din: boolean;
  signal op_mem_32_22_back: boolean;
  signal op_mem_32_22_push_front_pop_back_en: std_logic;
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  op_mem_32_22_back <= op_mem_32_22(0);
  proc_op_mem_32_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_32_22_push_front_pop_back_en = '1')) then
        op_mem_32_22(0) <= op_mem_32_22_front_din;
      end if;
    end if;
  end process proc_op_mem_32_22;
  result_12_3_rel <= a_1_31 = b_1_34;
  op_mem_32_22_front_din <= result_12_3_rel;
  op_mem_32_22_push_front_pop_back_en <= '1';
  op <= boolean_to_vector(op_mem_32_22_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_83ca2c6a3c is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_83ca2c6a3c;


architecture behavior of relational_83ca2c6a3c is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  type array_type_op_mem_32_22 is array (0 to (4 - 1)) of boolean;
  signal op_mem_32_22: array_type_op_mem_32_22 := (
    false,
    false,
    false,
    false);
  signal op_mem_32_22_front_din: boolean;
  signal op_mem_32_22_back: boolean;
  signal op_mem_32_22_push_front_pop_back_en: std_logic;
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  op_mem_32_22_back <= op_mem_32_22(3);
  proc_op_mem_32_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_32_22_push_front_pop_back_en = '1')) then
        for i in 3 downto 1 loop
          op_mem_32_22(i) <= op_mem_32_22(i-1);
        end loop;
        op_mem_32_22(0) <= op_mem_32_22_front_din;
      end if;
    end if;
  end process proc_op_mem_32_22;
  result_12_3_rel <= a_1_31 = b_1_34;
  op_mem_32_22_front_din <= result_12_3_rel;
  op_mem_32_22_push_front_pop_back_en <= '1';
  op <= boolean_to_vector(op_mem_32_22_back);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_2acadf5a08d72e0ee15ce4e1ac741dc6 is
  port(
    ce:in std_logic;
    ce_1400000:in std_logic;
    ce_2800000:in std_logic;
    ce_logic_1400000:in std_logic;
    clk:in std_logic;
    clk_1400000:in std_logic;
    clk_2800000:in std_logic;
    clk_logic_1400000:in std_logic;
    event_s_data_chanid_incorrect:out std_logic;
    m_axis_data_tdata:out std_logic_vector(24 downto 0);
    m_axis_data_tuser_chanid:out std_logic_vector(1 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    s_axis_data_tuser_chanid:in std_logic_vector(1 downto 0);
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_2acadf5a08d72e0ee15ce4e1ac741dc6;


architecture behavior of xlfir_compiler_2acadf5a08d72e0ee15ce4e1ac741dc6  is
  component fr_cmplr_v6_3_8e79a078fc118dc6
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_s_data_chanid_incorrect:out std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tuser:out std_logic_vector(1 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tuser:in std_logic_vector(1 downto 0);
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tuser_chanid_ps_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
signal s_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(24 downto 0);
  m_axis_data_tuser_chanid_ps_net <= m_axis_data_tuser_net(1 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata;
  s_axis_data_tuser_net(1 downto 0) <= s_axis_data_tuser_chanid;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_2800000,
        clr => '0',
        clk => clk_2800000,
        o => m_axis_data_tdata
    );
  m_axis_data_tuser_chanid_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 2,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chanid_ps_net,
        ce => ce_2800000,
        clr => '0',
        clk => clk_2800000,
        o => m_axis_data_tuser_chanid
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_2800000,
        clr => '0',
        clk => clk_2800000,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_2800000,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_8e79a078fc118dc6_instance : fr_cmplr_v6_3_8e79a078fc118dc6
    port map(
      aclk=>clk,
      aclken=>ce,
      event_s_data_chanid_incorrect=>event_s_data_chanid_incorrect,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tuser=>s_axis_data_tuser_net,
      s_axis_data_tvalid=>ce_logic_1400000
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlcic_compiler_6efc67831a277bdb0701519c5a976f20 is
  port(
    ce:in std_logic;
    ce_1400000:in std_logic;
    ce_560:in std_logic;
    ce_logic_560:in std_logic;
    clk:in std_logic;
    clk_1400000:in std_logic;
    clk_560:in std_logic;
    clk_logic_560:in std_logic;
    event_tlast_missing:out std_logic;
    event_tlast_unexpected:out std_logic;
    m_axis_data_tdata_data:out std_logic_vector(60 downto 0);
    m_axis_data_tlast:out std_logic;
    m_axis_data_tuser_chan_out:out std_logic_vector(1 downto 0);
    m_axis_data_tuser_chan_sync:out std_logic_vector(0 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_data:in std_logic_vector(23 downto 0);
    s_axis_data_tlast:in std_logic;
    s_axis_data_tready:out std_logic
  );
end xlcic_compiler_6efc67831a277bdb0701519c5a976f20;


architecture behavior of xlcic_compiler_6efc67831a277bdb0701519c5a976f20  is
  component cc_cmplr_v3_0_e58a4eb9f6488d2d
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_tlast_missing:out std_logic;
      event_tlast_unexpected:out std_logic;
      m_axis_data_tdata:out std_logic_vector(63 downto 0);
      m_axis_data_tlast:out std_logic;
      m_axis_data_tuser:out std_logic_vector(15 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tlast:in std_logic;
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net: std_logic_vector(60 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_captured: std_logic_vector(60 downto 0) := (others=>'0');
signal m_axis_data_tdata_data_ps_net_or_captured_net: std_logic_vector(60 downto 0) := (others=>'0');
signal m_axis_data_tlast_ps_net: std_logic := '0';
signal m_axis_data_tlast_ps_net_captured: std_logic := '0';
signal m_axis_data_tlast_ps_net_or_captured_net: std_logic := '0';
signal m_axis_data_tuser_net: std_logic_vector(15 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net_captured: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_sync_ps_net_or_captured_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net_captured: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tuser_chan_out_ps_net_or_captured_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_data_ps_net <= m_axis_data_tdata_net(60 downto 0);
  m_axis_data_tuser_chan_sync_ps_net <= m_axis_data_tuser_net(8 downto 8);
  m_axis_data_tuser_chan_out_ps_net <= m_axis_data_tuser_net(1 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_data;
  m_axis_data_tdata_data_ps_net_or_captured_net <= m_axis_data_tdata_data_ps_net or m_axis_data_tdata_data_ps_net_captured;
m_axis_data_tdata_data_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 61,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net_or_captured_net,
        ce => ce_1400000,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tdata_data
    );
m_axis_data_tdata_data_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 61,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_data_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tdata_data_ps_net_captured
    );
  m_axis_data_tlast_ps_net_or_captured_net <= m_axis_data_tlast_ps_net or m_axis_data_tlast_ps_net_captured;
m_axis_data_tlast_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tlast_ps_net_or_captured_net,
        ce => ce_1400000,
        clr => '0',
        clk => clk_1400000,
        o(0) => m_axis_data_tlast
    );
m_axis_data_tlast_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tlast_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1400000,
        o(0) => m_axis_data_tlast_ps_net_captured
    );
  m_axis_data_tuser_chan_sync_ps_net_or_captured_net <= m_axis_data_tuser_chan_sync_ps_net or m_axis_data_tuser_chan_sync_ps_net_captured;
m_axis_data_tuser_chan_sync_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_sync_ps_net_or_captured_net,
        ce => ce_1400000,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tuser_chan_sync
    );
m_axis_data_tuser_chan_sync_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_sync_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tuser_chan_sync_ps_net_captured
    );
  m_axis_data_tuser_chan_out_ps_net_or_captured_net <= m_axis_data_tuser_chan_out_ps_net or m_axis_data_tuser_chan_out_ps_net_captured;
m_axis_data_tuser_chan_out_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 2,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_out_ps_net_or_captured_net,
        ce => ce_1400000,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tuser_chan_out
    );
m_axis_data_tuser_chan_out_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 2,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chan_out_ps_net,
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1400000,
        o => m_axis_data_tuser_chan_out_ps_net_captured
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_1400000,
        clr => '0',
        clk => clk_1400000,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_1400000,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  cc_cmplr_v3_0_e58a4eb9f6488d2d_instance : cc_cmplr_v3_0_e58a4eb9f6488d2d
    port map(
      aclk=>clk,
      aclken=>ce,
      event_tlast_missing=>event_tlast_missing,
      event_tlast_unexpected=>event_tlast_unexpected,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tlast=>m_axis_data_tlast_ps_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tlast=>s_axis_data_tlast,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>ce_logic_560
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_1da691037bdf8c1b85b3b4502d6e9610 is
  port(
    ce:in std_logic;
    ce_2800000:in std_logic;
    ce_5600000:in std_logic;
    ce_logic_2800000:in std_logic;
    clk:in std_logic;
    clk_2800000:in std_logic;
    clk_5600000:in std_logic;
    clk_logic_2800000:in std_logic;
    event_s_data_chanid_incorrect:out std_logic;
    m_axis_data_tdata:out std_logic_vector(24 downto 0);
    m_axis_data_tuser_chanid:out std_logic_vector(1 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    s_axis_data_tuser_chanid:in std_logic_vector(1 downto 0);
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_1da691037bdf8c1b85b3b4502d6e9610;


architecture behavior of xlfir_compiler_1da691037bdf8c1b85b3b4502d6e9610  is
  component fr_cmplr_v6_3_15ffe94f3ff4129f
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_s_data_chanid_incorrect:out std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tuser:out std_logic_vector(1 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(23 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tuser:in std_logic_vector(1 downto 0);
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tuser_chanid_ps_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(23 downto 0) := (others=>'0');
signal s_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(24 downto 0);
  m_axis_data_tuser_chanid_ps_net <= m_axis_data_tuser_net(1 downto 0);
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata;
  s_axis_data_tuser_net(1 downto 0) <= s_axis_data_tuser_chanid;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_5600000,
        clr => '0',
        clk => clk_5600000,
        o => m_axis_data_tdata
    );
  m_axis_data_tuser_chanid_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 2,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chanid_ps_net,
        ce => ce_5600000,
        clr => '0',
        clk => clk_5600000,
        o => m_axis_data_tuser_chanid
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_5600000,
        clr => '0',
        clk => clk_5600000,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_5600000,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_15ffe94f3ff4129f_instance : fr_cmplr_v6_3_15ffe94f3ff4129f
    port map(
      aclk=>clk,
      aclken=>ce,
      event_s_data_chanid_incorrect=>event_s_data_chanid_incorrect,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tuser=>s_axis_data_tuser_net,
      s_axis_data_tvalid=>ce_logic_2800000
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_f7093b59b74f3d511e09195b077ec73c is
  port(
    ce:in std_logic;
    ce_35:in std_logic;
    ce_logic_1:in std_logic;
    clk:in std_logic;
    clk_35:in std_logic;
    clk_logic_1:in std_logic;
    event_s_data_chanid_incorrect:out std_logic;
    m_axis_data_tdata_path0:out std_logic_vector(24 downto 0);
    m_axis_data_tdata_path1:out std_logic_vector(24 downto 0);
    m_axis_data_tuser_chanid:out std_logic_vector(0 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata_path0:in std_logic_vector(23 downto 0);
    s_axis_data_tdata_path1:in std_logic_vector(23 downto 0);
    s_axis_data_tready:out std_logic;
    s_axis_data_tuser_chanid:in std_logic_vector(0 downto 0);
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_f7093b59b74f3d511e09195b077ec73c;


architecture behavior of xlfir_compiler_f7093b59b74f3d511e09195b077ec73c  is
  component fr_cmplr_v6_3_2b018066c9a0cd8a
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_s_data_chanid_incorrect:out std_logic;
      m_axis_data_tdata:out std_logic_vector(63 downto 0);
      m_axis_data_tuser:out std_logic_vector(0 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(47 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tuser:in std_logic_vector(0 downto 0);
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(63 downto 0) := (others=>'0');
signal m_axis_data_tdata_path1_ps_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tdata_path0_ps_net: std_logic_vector(24 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tuser_chanid_ps_net: std_logic_vector(0 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(47 downto 0) := (others=>'0');
signal s_axis_data_tuser_net: std_logic_vector(0 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_path1_ps_net <= m_axis_data_tdata_net(56 downto 32);
  m_axis_data_tdata_path0_ps_net <= m_axis_data_tdata_net(24 downto 0);
  m_axis_data_tuser_chanid_ps_net <= m_axis_data_tuser_net(0 downto 0);
  s_axis_data_tdata_net(47 downto 24) <= s_axis_data_tdata_path1;
  s_axis_data_tdata_net(23 downto 0) <= s_axis_data_tdata_path0;
  s_axis_data_tuser_net(0 downto 0) <= s_axis_data_tuser_chanid;
  m_axis_data_tdata_path1_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_path1_ps_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35,
        o => m_axis_data_tdata_path1
    );
  m_axis_data_tdata_path0_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 25,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_path0_ps_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35,
        o => m_axis_data_tdata_path0
    );
  m_axis_data_tuser_chanid_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chanid_ps_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35,
        o => m_axis_data_tuser_chanid
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_35,
        clr => '0',
        clk => clk_35,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_35,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_2b018066c9a0cd8a_instance : fr_cmplr_v6_3_2b018066c9a0cd8a
    port map(
      aclk=>clk,
      aclken=>ce,
      event_s_data_chanid_incorrect=>event_s_data_chanid_incorrect,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tuser=>s_axis_data_tuser_net,
      s_axis_data_tvalid=>ce_logic_1
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f062741975 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((24 - 1) downto 0);
    d1 : in std_logic_vector((24 - 1) downto 0);
    d2 : in std_logic_vector((24 - 1) downto 0);
    d3 : in std_logic_vector((24 - 1) downto 0);
    y : out std_logic_vector((24 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f062741975;


architecture behavior of mux_f062741975 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((24 - 1) downto 0);
  signal d1_1_27: std_logic_vector((24 - 1) downto 0);
  signal d2_1_30: std_logic_vector((24 - 1) downto 0);
  signal d3_1_33: std_logic_vector((24 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((24 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlcounter_free is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free ;
architecture behavior of xlcounter_free is
  component cntr_11_0_eb46eda57512a5a4
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of cntr_11_0_eb46eda57512a5a4:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_eb46eda57512a5a4:
    component is "true";
  attribute box_type of cntr_11_0_eb46eda57512a5a4:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_eb46eda57512a5a4")) generate
    core_instance0: cntr_11_0_eb46eda57512a5a4
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_187c900130 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((26 - 1) downto 0);
    d1 : in std_logic_vector((26 - 1) downto 0);
    d2 : in std_logic_vector((26 - 1) downto 0);
    d3 : in std_logic_vector((26 - 1) downto 0);
    y : out std_logic_vector((26 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_187c900130;


architecture behavior of mux_187c900130 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((26 - 1) downto 0);
  signal d1_1_27: std_logic_vector((26 - 1) downto 0);
  signal d2_1_30: std_logic_vector((26 - 1) downto 0);
  signal d3_1_33: std_logic_vector((26 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((26 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_60ea556961 is
  port (
    input_port : in std_logic_vector((25 - 1) downto 0);
    output_port : out std_logic_vector((25 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_60ea556961;


architecture behavior of reinterpret_60ea556961 is
  signal input_port_1_40: unsigned((25 - 1) downto 0);
  signal output_port_5_5_force: signed((25 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity bitbasher_a756ba0096 is
  port (
    din : in std_logic_vector((26 - 1) downto 0);
    dout : out std_logic_vector((25 - 1) downto 0);
    vld_out : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end bitbasher_a756ba0096;


architecture behavior of bitbasher_a756ba0096 is
  signal din_1_37: unsigned((26 - 1) downto 0);
  signal slice_5_31: unsigned((25 - 1) downto 0);
  signal fulldout_5_1_concat: unsigned((25 - 1) downto 0);
  signal slice_6_44: unsigned((1 - 1) downto 0);
  signal concat_6_35: unsigned((1 - 1) downto 0);
  signal fullvld_out_6_1_concat: unsigned((1 - 1) downto 0);
begin
  din_1_37 <= std_logic_vector_to_unsigned(din);
  slice_5_31 <= u2u_slice(din_1_37, 24, 0);
  fulldout_5_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(slice_5_31));
  slice_6_44 <= u2u_slice(din_1_37, 25, 25);
  concat_6_35 <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(slice_6_44));
  fullvld_out_6_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(concat_6_35));
  dout <= unsigned_to_std_logic_vector(fulldout_5_1_concat);
  vld_out <= unsigned_to_std_logic_vector(fullvld_out_6_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_80f90b97d0 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_80f90b97d0;


architecture behavior of logical_80f90b97d0 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlpassthrough is
    generic (
        din_width    : integer := 16;
        dout_width   : integer := 16
        );
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlpassthrough;
architecture passthrough_arch of xlpassthrough is
begin
  dout <= din;
end passthrough_arch;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity expr_375d7bbece is
  port (
    a : in std_logic_vector((1 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    c : in std_logic_vector((1 - 1) downto 0);
    dout : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end expr_375d7bbece;


architecture behavior of expr_375d7bbece is
  signal a_1_24: boolean;
  signal b_1_27: boolean;
  signal c_1_30: boolean;
  signal bit_6_36: boolean;
  signal fulldout_6_2_bit: boolean;
begin
  a_1_24 <= ((a) = "1");
  b_1_27 <= ((b) = "1");
  c_1_30 <= ((c) = "1");
  bit_6_36 <= ((boolean_to_vector(b_1_27) and boolean_to_vector(a_1_24)) = "1");
  fulldout_6_2_bit <= ((boolean_to_vector(c_1_30) and boolean_to_vector(bit_6_36)) = "1");
  dout <= boolean_to_vector(fulldout_6_2_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc is
  port(
    ce:in std_logic;
    clk:in std_logic;
    m_axis_dout_tdata_fractional:out std_logic_vector(24 downto 0);
    m_axis_dout_tdata_quotient:out std_logic_vector(25 downto 0);
    m_axis_dout_tvalid:out std_logic;
    s_axis_dividend_tdata_dividend:in std_logic_vector(25 downto 0);
    s_axis_dividend_tready:out std_logic;
    s_axis_dividend_tvalid:in std_logic;
    s_axis_divisor_tdata_divisor:in std_logic_vector(25 downto 0);
    s_axis_divisor_tready:out std_logic;
    s_axis_divisor_tvalid:in std_logic
  );
end xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc;


architecture behavior of xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc  is
  component dv_gn_v4_0_dc31160d1288a80d
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      m_axis_dout_tdata:out std_logic_vector(55 downto 0);
      m_axis_dout_tvalid:out std_logic;
      s_axis_dividend_tdata:in std_logic_vector(31 downto 0);
      s_axis_dividend_tready:out std_logic;
      s_axis_dividend_tvalid:in std_logic;
      s_axis_divisor_tdata:in std_logic_vector(31 downto 0);
      s_axis_divisor_tready:out std_logic;
      s_axis_divisor_tvalid:in std_logic
    );
end component;
signal m_axis_dout_tdata_net: std_logic_vector(55 downto 0) := (others=>'0');
signal s_axis_dividend_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal s_axis_divisor_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  m_axis_dout_tdata_quotient <= m_axis_dout_tdata_net(50 downto 25);
  m_axis_dout_tdata_fractional <= m_axis_dout_tdata_net(24 downto 0);
  s_axis_dividend_tdata_net(25 downto 0) <= s_axis_dividend_tdata_dividend;
  s_axis_divisor_tdata_net(25 downto 0) <= s_axis_divisor_tdata_divisor;
  dv_gn_v4_0_dc31160d1288a80d_instance : dv_gn_v4_0_dc31160d1288a80d
    port map(
      aclk=>clk,
      aclken=>ce,
      m_axis_dout_tdata=>m_axis_dout_tdata_net,
      m_axis_dout_tvalid=>m_axis_dout_tvalid,
      s_axis_dividend_tdata=>s_axis_dividend_tdata_net,
      s_axis_dividend_tready=>s_axis_dividend_tready,
      s_axis_dividend_tvalid=>s_axis_dividend_tvalid,
      s_axis_divisor_tdata=>s_axis_divisor_tdata_net,
      s_axis_divisor_tready=>s_axis_divisor_tready,
      s_axis_divisor_tvalid=>s_axis_divisor_tvalid
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_040ef1b598 is
  port (
    input_port : in std_logic_vector((26 - 1) downto 0);
    output_port : out std_logic_vector((26 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_040ef1b598;


architecture behavior of reinterpret_040ef1b598 is
  signal input_port_1_40: signed((26 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port <= signed_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_416cfcae1e is
  port (
    a : in std_logic_vector((26 - 1) downto 0);
    b : in std_logic_vector((26 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_416cfcae1e;


architecture behavior of relational_416cfcae1e is
  signal a_1_31: signed((26 - 1) downto 0);
  signal b_1_34: signed((26 - 1) downto 0);
  type array_type_op_mem_32_22 is array (0 to (1 - 1)) of boolean;
  signal op_mem_32_22: array_type_op_mem_32_22 := (
    0 => false);
  signal op_mem_32_22_front_din: boolean;
  signal op_mem_32_22_back: boolean;
  signal op_mem_32_22_push_front_pop_back_en: std_logic;
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_signed(a);
  b_1_34 <= std_logic_vector_to_signed(b);
  op_mem_32_22_back <= op_mem_32_22(0);
  proc_op_mem_32_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_32_22_push_front_pop_back_en = '1')) then
        op_mem_32_22(0) <= op_mem_32_22_front_din;
      end if;
    end if;
  end process proc_op_mem_32_22;
  result_18_3_rel <= a_1_31 > b_1_34;
  op_mem_32_22_front_din <= result_18_3_rel;
  op_mem_32_22_push_front_pop_back_en <= '1';
  op <= boolean_to_vector(op_mem_32_22_back);
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.4 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub;
architecture behavior of xladdsub is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_293aa5f110d040c2
    port (
          a: in std_logic_vector(25 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(25 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_293aa5f110d040c2:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_293aa5f110d040c2:
    component is "true";
  attribute box_type of addsb_11_0_293aa5f110d040c2:
    component  is "black_box";
  component addsb_11_0_44053abf11139d96
    port (
          a: in std_logic_vector(26 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(26 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_44053abf11139d96:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_44053abf11139d96:
    component is "true";
  attribute box_type of addsb_11_0_44053abf11139d96:
    component  is "black_box";
  component addsb_11_0_3537d66a2361cd1e
    port (
          a: in std_logic_vector(26 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(26 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_3537d66a2361cd1e:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_3537d66a2361cd1e:
    component is "true";
  attribute box_type of addsb_11_0_3537d66a2361cd1e:
    component  is "black_box";
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_293aa5f110d040c2")) generate
    core_instance0: addsb_11_0_293aa5f110d040c2
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp1: if ((core_name0 = "addsb_11_0_44053abf11139d96")) generate
    core_instance1: addsb_11_0_44053abf11139d96
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_3537d66a2361cd1e")) generate
    core_instance2: addsb_11_0_3537d66a2361cd1e
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_43e7f055fa is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((25 - 1) downto 0);
    y : out std_logic_vector((26 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_43e7f055fa;


architecture behavior of concat_43e7f055fa is
  signal in0_1_23: boolean;
  signal in1_1_27: unsigned((25 - 1) downto 0);
  signal y_2_1_concat: unsigned((26 - 1) downto 0);
begin
  in0_1_23 <= ((in0) = "1");
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(boolean_to_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_c3c0e847be is
  port (
    input_port : in std_logic_vector((25 - 1) downto 0);
    output_port : out std_logic_vector((25 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_c3c0e847be;


architecture behavior of reinterpret_c3c0e847be is
  signal input_port_1_40: signed((25 - 1) downto 0);
  signal output_port_5_5_force: unsigned((25 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfir_compiler_eebfed0cb0075aa32aca169bb967f58b is
  port(
    ce:in std_logic;
    ce_5600000:in std_logic;
    ce_56000000:in std_logic;
    ce_logic_5600000:in std_logic;
    clk:in std_logic;
    clk_5600000:in std_logic;
    clk_56000000:in std_logic;
    clk_logic_5600000:in std_logic;
    event_s_data_chanid_incorrect:out std_logic;
    m_axis_data_tdata:out std_logic_vector(25 downto 0);
    m_axis_data_tuser_chanid:out std_logic_vector(1 downto 0);
    m_axis_data_tvalid:out std_logic;
    s_axis_data_tdata:in std_logic_vector(24 downto 0);
    s_axis_data_tready:out std_logic;
    s_axis_data_tuser_chanid:in std_logic_vector(1 downto 0);
    src_ce:in std_logic;
    src_clk:in std_logic
  );
end xlfir_compiler_eebfed0cb0075aa32aca169bb967f58b;


architecture behavior of xlfir_compiler_eebfed0cb0075aa32aca169bb967f58b  is
  component fr_cmplr_v6_3_b1697e0c92d2e32a
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      event_s_data_chanid_incorrect:out std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tuser:out std_logic_vector(1 downto 0);
      m_axis_data_tvalid:out std_logic;
      s_axis_data_tdata:in std_logic_vector(31 downto 0);
      s_axis_data_tready:out std_logic;
      s_axis_data_tuser:in std_logic_vector(1 downto 0);
      s_axis_data_tvalid:in std_logic
    );
end component;
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tdata_ps_net: std_logic_vector(25 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tuser_chanid_ps_net: std_logic_vector(1 downto 0) := (others=>'0');
signal m_axis_data_tvalid_ps_net: std_logic := '0';
signal m_axis_data_tvalid_ps_net_captured: std_logic := '0';
signal m_axis_data_tvalid_ps_net_or_captured_net: std_logic := '0';
signal s_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal s_axis_data_tuser_net: std_logic_vector(1 downto 0) := (others=>'0');
begin
  m_axis_data_tdata_ps_net <= m_axis_data_tdata_net(25 downto 0);
  m_axis_data_tuser_chanid_ps_net <= m_axis_data_tuser_net(1 downto 0);
  s_axis_data_tdata_net(24 downto 0) <= s_axis_data_tdata;
  s_axis_data_tuser_net(1 downto 0) <= s_axis_data_tuser_chanid;
  m_axis_data_tdata_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 26,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tdata_ps_net,
        ce => ce_56000000,
        clr => '0',
        clk => clk_56000000,
        o => m_axis_data_tdata
    );
  m_axis_data_tuser_chanid_ps_net_synchronizer : entity work.synth_reg_w_init
    generic map(
        width => 2,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i => m_axis_data_tuser_chanid_ps_net,
        ce => ce_56000000,
        clr => '0',
        clk => clk_56000000,
        o => m_axis_data_tuser_chanid
    );
  m_axis_data_tvalid_ps_net_or_captured_net <= m_axis_data_tvalid_ps_net or m_axis_data_tvalid_ps_net_captured;
m_axis_data_tvalid_ps_net_synchronizer_1 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => m_axis_data_tvalid_ps_net_or_captured_net,
        ce => ce_56000000,
        clr => '0',
        clk => clk_56000000,
        o(0) => m_axis_data_tvalid
    );
m_axis_data_tvalid_ps_net_synchronizer_2 : entity work.synth_reg_w_init
    generic map(
        width => 1,
        init_index => 0,
        init_value => "0",
        latency => 1
    )
    port map (
        i(0) => '1',
        ce => m_axis_data_tvalid_ps_net,
        clr => '0',
        clk => clk_56000000,
        o(0) => m_axis_data_tvalid_ps_net_captured
    );
  fr_cmplr_v6_3_b1697e0c92d2e32a_instance : fr_cmplr_v6_3_b1697e0c92d2e32a
    port map(
      aclk=>clk,
      aclken=>ce,
      event_s_data_chanid_incorrect=>event_s_data_chanid_incorrect,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid_ps_net,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tuser=>s_axis_data_tuser_net,
      s_axis_data_tvalid=>ce_logic_5600000
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/BPF/zero_filling1"

entity zero_filling1_entity_d0ac9899b1 is
  port (
    in1: in std_logic_vector(15 downto 0);
    out1: out std_logic_vector(23 downto 0)
  );
end zero_filling1_entity_d0ac9899b1;

architecture structural of zero_filling1_entity_d0ac9899b1 is
  signal concat_y_net: std_logic_vector(23 downto 0);
  signal constant_op_net: std_logic_vector(7 downto 0);
  signal register1_q_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(7 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  register1_q_net_x0 <= in1;
  out1 <= reinterpret2_output_port_net_x0;

  concat: entity work.concat_cd3162dc0d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net
    );

  constant_x0: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  reinterpret: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => register1_q_net_x0,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_f21e7f2ddf
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => constant_op_net,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_4bf1ad328a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => concat_y_net,
      output_port => reinterpret2_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/BPF"

entity bpf_entity_d31c4af409 is
  port (
    din_ch0: in std_logic_vector(15 downto 0);
    din_ch1: in std_logic_vector(15 downto 0);
    din_ch2: in std_logic_vector(15 downto 0);
    din_ch3: in std_logic_vector(15 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0);
    dout_ch2: out std_logic_vector(23 downto 0);
    dout_ch3: out std_logic_vector(23 downto 0)
  );
end bpf_entity_d31c4af409;

architecture structural of bpf_entity_d31c4af409 is
  signal register1_q_net_x1: std_logic_vector(15 downto 0);
  signal register2_q_net_x1: std_logic_vector(15 downto 0);
  signal register3_q_net_x1: std_logic_vector(15 downto 0);
  signal register_q_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x4: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x5: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x6: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x7: std_logic_vector(23 downto 0);

begin
  register_q_net_x1 <= din_ch0;
  register1_q_net_x1 <= din_ch1;
  register2_q_net_x1 <= din_ch2;
  register3_q_net_x1 <= din_ch3;
  dout_ch0 <= reinterpret2_output_port_net_x7;
  dout_ch1 <= reinterpret2_output_port_net_x4;
  dout_ch2 <= reinterpret2_output_port_net_x5;
  dout_ch3 <= reinterpret2_output_port_net_x6;

  zero_filling1_d0ac9899b1: entity work.zero_filling1_entity_d0ac9899b1
    port map (
      in1 => register1_q_net_x1,
      out1 => reinterpret2_output_port_net_x4
    );

  zero_filling2_d7e27e9bae: entity work.zero_filling1_entity_d0ac9899b1
    port map (
      in1 => register2_q_net_x1,
      out1 => reinterpret2_output_port_net_x5
    );

  zero_filling3_1ae3b6c91e: entity work.zero_filling1_entity_d0ac9899b1
    port map (
      in1 => register3_q_net_x1,
      out1 => reinterpret2_output_port_net_x6
    );

  zero_filling4_6d7b2d0c57: entity work.zero_filling1_entity_d0ac9899b1
    port map (
      in1 => register_q_net_x1,
      out1 => reinterpret2_output_port_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/DDS_sub/TDM_dds_ch01_cosine"

entity tdm_dds_ch01_cosine_entity_4b8bfc9243 is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_logic_1: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    din_ch0: in std_logic_vector(23 downto 0);
    rst: in std_logic;
    dout: out std_logic_vector(23 downto 0)
  );
end tdm_dds_ch01_cosine_entity_4b8bfc9243;

architecture structural of tdm_dds_ch01_cosine_entity_4b8bfc9243 is
  signal black_box_cos_o_net_x0: std_logic_vector(23 downto 0);
  signal ce_1_sg_x0: std_logic;
  signal ce_2_sg_x0: std_logic;
  signal ce_logic_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal clk_2_sg_x0: std_logic;
  signal clock_enable_probe_q_net: std_logic;
  signal constant11_op_net_x0: std_logic;
  signal mux_sel1_op_net: std_logic;
  signal mux_y_net: std_logic_vector(23 downto 0);
  signal register2_q_net: std_logic_vector(23 downto 0);
  signal register3_q_net: std_logic_vector(23 downto 0);
  signal register4_q_net: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal up_sample_ch0_q_net: std_logic_vector(23 downto 0);
  signal up_sample_ch1_q_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  ce_2_sg_x0 <= ce_2;
  ce_logic_1_sg_x0 <= ce_logic_1;
  clk_1_sg_x0 <= clk_1;
  clk_2_sg_x0 <= clk_2;
  black_box_cos_o_net_x0 <= din_ch0;
  constant11_op_net_x0 <= rst;
  dout <= register_q_net_x0;

  clock_enable_probe: entity work.xlceprobe
    generic map (
      d_width => 24,
      q_width => 1
    )
    port map (
      ce => ce_logic_1_sg_x0,
      clk => clk_1_sg_x0,
      d => register2_q_net,
      q(0) => clock_enable_probe_q_net
    );

  mux: entity work.mux_a2121d82da
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register2_q_net,
      d1 => register3_q_net,
      sel(0) => register4_q_net,
      y => mux_y_net
    );

  mux_sel1: entity work.counter_41314d726b
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => clock_enable_probe_q_net,
      rst(0) => constant11_op_net_x0,
      op(0) => mux_sel1_op_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => up_sample_ch0_q_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => up_sample_ch1_q_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => mux_sel1_op_net,
      en => "1",
      rst => "0",
      q(0) => register4_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => mux_y_net,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

  up_sample_ch0: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => black_box_cos_o_net_x0,
      dest_ce => ce_1_sg_x0,
      dest_clk => clk_1_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x0,
      src_clk => clk_2_sg_x0,
      src_clr => '0',
      q => up_sample_ch0_q_net
    );

  up_sample_ch1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => black_box_cos_o_net_x0,
      dest_ce => ce_1_sg_x0,
      dest_clk => clk_1_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x0,
      src_clk => clk_2_sg_x0,
      src_clr => '0',
      q => up_sample_ch1_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
use work.dsp_cores_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/DDS_sub"

entity dds_sub_entity_a4b6b880f6 is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_logic_1: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    dds_01_cosine: out std_logic_vector(23 downto 0);
    dds_01_sine: out std_logic_vector(23 downto 0);
    dds_23_cosine: out std_logic_vector(23 downto 0);
    dds_23_sine: out std_logic_vector(23 downto 0)
  );
end dds_sub_entity_a4b6b880f6;

architecture structural of dds_sub_entity_a4b6b880f6 is
  signal black_box_cos_o_net_x1: std_logic_vector(23 downto 0);
  signal black_box_sin_o_net_x1: std_logic_vector(23 downto 0);
  signal ce_1_sg_x4: std_logic;
  signal ce_2_sg_x4: std_logic;
  signal ce_logic_1_sg_x4: std_logic;
  signal clk_1_sg_x4: std_logic;
  signal clk_2_sg_x4: std_logic;
  signal constant11_op_net_x0: std_logic;
  signal constant16_op_net_x0: std_logic;
  signal constant17_op_net_x0: std_logic;
  signal constant3_op_net: std_logic;
  signal constant7_op_net_x0: std_logic;
  signal register_q_net_x4: std_logic_vector(23 downto 0);
  signal register_q_net_x5: std_logic_vector(23 downto 0);
  signal register_q_net_x6: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x4 <= ce_1;
  ce_2_sg_x4 <= ce_2;
  ce_logic_1_sg_x4 <= ce_logic_1;
  clk_1_sg_x4 <= clk_1;
  clk_2_sg_x4 <= clk_2;
  dds_01_cosine <= register_q_net_x4;
  dds_01_sine <= register_q_net_x5;
  dds_23_cosine <= register_q_net_x6;
  dds_23_sine <= register_q_net_x7;

  black_box: entity work.fixed_dds
    generic map (
      g_cos_file => f_dds_cos_file(c_machine_name),
      g_dither => false,
      g_number_of_points => f_dds_num_points(c_machine_name),
      g_output_width => 24,
      g_sin_file => f_dds_sin_file(c_machine_name)
    )
    port map (
      ce_i => ce_2_sg_x4,
      clk_i => clk_2_sg_x4,
      rst_n_i => constant3_op_net,
      cos_o => black_box_cos_o_net_x1,
      sin_o => black_box_sin_o_net_x1
    );

  constant11: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant11_op_net_x0
    );

  constant16: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant16_op_net_x0
    );

  constant17: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant17_op_net_x0
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant7: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant7_op_net_x0
    );

  tdm_dds_ch01_cosine_4b8bfc9243: entity work.tdm_dds_ch01_cosine_entity_4b8bfc9243
    port map (
      ce_1 => ce_1_sg_x4,
      ce_2 => ce_2_sg_x4,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x4,
      clk_2 => clk_2_sg_x4,
      din_ch0 => black_box_cos_o_net_x1,
      rst => constant11_op_net_x0,
      dout => register_q_net_x4
    );

  tdm_dds_ch01_sine_1129eb9762: entity work.tdm_dds_ch01_cosine_entity_4b8bfc9243
    port map (
      ce_1 => ce_1_sg_x4,
      ce_2 => ce_2_sg_x4,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x4,
      clk_2 => clk_2_sg_x4,
      din_ch0 => black_box_sin_o_net_x1,
      rst => constant7_op_net_x0,
      dout => register_q_net_x5
    );

  tdm_dds_ch23_cosine_398d5cee32: entity work.tdm_dds_ch01_cosine_entity_4b8bfc9243
    port map (
      ce_1 => ce_1_sg_x4,
      ce_2 => ce_2_sg_x4,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x4,
      clk_2 => clk_2_sg_x4,
      din_ch0 => black_box_cos_o_net_x1,
      rst => constant16_op_net_x0,
      dout => register_q_net_x6
    );

  tdm_dds_ch23_sine_782ff6a42a: entity work.tdm_dds_ch01_cosine_entity_4b8bfc9243
    port map (
      ce_1 => ce_1_sg_x4,
      ce_2 => ce_2_sg_x4,
      ce_logic_1 => ce_logic_1_sg_x4,
      clk_1 => clk_1_sg_x4,
      clk_2 => clk_2_sg_x4,
      din_ch0 => black_box_sin_o_net_x1,
      rst => constant17_op_net_x0,
      dout => register_q_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/TDDM_fofb_amp_4ch/TDDM_fofb_amp0"

entity tddm_fofb_amp0_entity_fd74c6ad6e is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ch_in: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_fofb_amp0_entity_fd74c6ad6e;

architecture structural of tddm_fofb_amp0_entity_fd74c6ad6e is
  signal ce_1120_sg_x0: std_logic;
  signal ce_2240_sg_x0: std_logic;
  signal clk_1120_sg_x0: std_logic;
  signal clk_2240_sg_x0: std_logic;
  signal constant1_op_net: std_logic;
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register5_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1120_sg_x0 <= ce_1120;
  ce_2240_sg_x0 <= ce_2240;
  register1_q_net_x1 <= ch_in;
  clk_1120_sg_x0 <= clk_1120;
  clk_2240_sg_x0 <= clk_2240;
  register5_q_net_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_2240_sg_x0,
      dest_clk => clk_2240_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1120_sg_x0,
      src_clk => clk_1120_sg_x0,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_2240_sg_x0,
      dest_clk => clk_2240_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1120_sg_x0,
      src_clk => clk_1120_sg_x0,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x0,
      clk => clk_1120_sg_x0,
      d => register5_q_net_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x0,
      clk => clk_1120_sg_x0,
      d => register5_q_net_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => register1_q_net_x1,
      b(0) => constant_op_net,
      ce => ce_1120_sg_x0,
      clk => clk_1120_sg_x0,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_a892e1bf40
    port map (
      a(0) => register1_q_net_x1,
      b(0) => constant1_op_net,
      ce => ce_1120_sg_x0,
      clk => clk_1120_sg_x0,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/TDDM_fofb_amp_4ch"

entity tddm_fofb_amp_4ch_entity_2cc521a83f is
  port (
    amp_in0: in std_logic_vector(23 downto 0);
    amp_in1: in std_logic_vector(23 downto 0);
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ch_in0: in std_logic;
    ch_in1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    amp_out0: out std_logic_vector(23 downto 0);
    amp_out1: out std_logic_vector(23 downto 0);
    amp_out2: out std_logic_vector(23 downto 0);
    amp_out3: out std_logic_vector(23 downto 0)
  );
end tddm_fofb_amp_4ch_entity_2cc521a83f;

architecture structural of tddm_fofb_amp_4ch_entity_2cc521a83f is
  signal ce_1120_sg_x2: std_logic;
  signal ce_2240_sg_x2: std_logic;
  signal clk_1120_sg_x2: std_logic;
  signal clk_2240_sg_x2: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x4: std_logic;
  signal register5_q_net_x2: std_logic_vector(23 downto 0);
  signal register5_q_net_x3: std_logic_vector(23 downto 0);

begin
  register5_q_net_x2 <= amp_in0;
  register5_q_net_x3 <= amp_in1;
  ce_1120_sg_x2 <= ce_1120;
  ce_2240_sg_x2 <= ce_2240;
  register1_q_net_x3 <= ch_in0;
  register1_q_net_x4 <= ch_in1;
  clk_1120_sg_x2 <= clk_1120;
  clk_2240_sg_x2 <= clk_2240;
  amp_out0 <= down_sample2_q_net_x2;
  amp_out1 <= down_sample1_q_net_x2;
  amp_out2 <= down_sample2_q_net_x3;
  amp_out3 <= down_sample1_q_net_x3;

  tddm_fofb_amp0_fd74c6ad6e: entity work.tddm_fofb_amp0_entity_fd74c6ad6e
    port map (
      ce_1120 => ce_1120_sg_x2,
      ce_2240 => ce_2240_sg_x2,
      ch_in => register1_q_net_x3,
      clk_1120 => clk_1120_sg_x2,
      clk_2240 => clk_2240_sg_x2,
      din => register5_q_net_x2,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_fofb_amp1_61cbc8ec65: entity work.tddm_fofb_amp0_entity_fd74c6ad6e
    port map (
      ce_1120 => ce_1120_sg_x2,
      ce_2240 => ce_2240_sg_x2,
      ch_in => register1_q_net_x4,
      clk_1120 => clk_1120_sg_x2,
      clk_2240 => clk_2240_sg_x2,
      din => register5_q_net_x3,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_CORDIC/TDDM_tbt_cordic0/TDDM_tbt_cordic1"

entity tddm_tbt_cordic1_entity_b60a69fd9b is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ch_in: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic1_entity_b60a69fd9b;

architecture structural of tddm_tbt_cordic1_entity_b60a69fd9b is
  signal ce_1120_sg_x4: std_logic;
  signal ce_2240_sg_x4: std_logic;
  signal clk_1120_sg_x4: std_logic;
  signal clk_2240_sg_x4: std_logic;
  signal constant1_op_net: std_logic;
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register1_q_net_x5: std_logic;
  signal register4_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1120_sg_x4 <= ce_1120;
  ce_2240_sg_x4 <= ce_2240;
  register1_q_net_x5 <= ch_in;
  clk_1120_sg_x4 <= clk_1120;
  clk_2240_sg_x4 <= clk_2240;
  register4_q_net_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_2240_sg_x4,
      dest_clk => clk_2240_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1120_sg_x4,
      src_clk => clk_1120_sg_x4,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_2240_sg_x4,
      dest_clk => clk_2240_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1120_sg_x4,
      src_clk => clk_1120_sg_x4,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x4,
      clk => clk_1120_sg_x4,
      d => register4_q_net_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x4,
      clk => clk_1120_sg_x4,
      d => register4_q_net_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => register1_q_net_x5,
      b(0) => constant_op_net,
      ce => ce_1120_sg_x4,
      clk => clk_1120_sg_x4,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_a892e1bf40
    port map (
      a(0) => register1_q_net_x5,
      b(0) => constant1_op_net,
      ce => ce_1120_sg_x4,
      clk => clk_1120_sg_x4,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_CORDIC/TDDM_tbt_cordic0"

entity tddm_tbt_cordic0_entity_38de3613fe is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    fofb_cordic_ch_in: in std_logic;
    fofb_cordic_din: in std_logic_vector(23 downto 0);
    fofb_cordic_pin: in std_logic_vector(23 downto 0);
    fofb_cordic_data0_out: out std_logic_vector(23 downto 0);
    fofb_cordic_data1_out: out std_logic_vector(23 downto 0);
    fofb_cordic_phase0_out: out std_logic_vector(23 downto 0);
    fofb_cordic_phase1_out: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic0_entity_38de3613fe;

architecture structural of tddm_tbt_cordic0_entity_38de3613fe is
  signal ce_1120_sg_x5: std_logic;
  signal ce_2240_sg_x5: std_logic;
  signal clk_1120_sg_x5: std_logic;
  signal clk_2240_sg_x5: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal register1_q_net_x6: std_logic;
  signal register4_q_net_x1: std_logic_vector(23 downto 0);
  signal register5_q_net_x4: std_logic_vector(23 downto 0);

begin
  ce_1120_sg_x5 <= ce_1120;
  ce_2240_sg_x5 <= ce_2240;
  clk_1120_sg_x5 <= clk_1120;
  clk_2240_sg_x5 <= clk_2240;
  register1_q_net_x6 <= fofb_cordic_ch_in;
  register5_q_net_x4 <= fofb_cordic_din;
  register4_q_net_x1 <= fofb_cordic_pin;
  fofb_cordic_data0_out <= down_sample2_q_net_x2;
  fofb_cordic_data1_out <= down_sample1_q_net_x2;
  fofb_cordic_phase0_out <= down_sample2_q_net_x3;
  fofb_cordic_phase1_out <= down_sample1_q_net_x3;

  tddm_fofb_cordic0_int_516d0c2a22: entity work.tddm_fofb_amp0_entity_fd74c6ad6e
    port map (
      ce_1120 => ce_1120_sg_x5,
      ce_2240 => ce_2240_sg_x5,
      ch_in => register1_q_net_x6,
      clk_1120 => clk_1120_sg_x5,
      clk_2240 => clk_2240_sg_x5,
      din => register5_q_net_x4,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_tbt_cordic1_b60a69fd9b: entity work.tddm_tbt_cordic1_entity_b60a69fd9b
    port map (
      ce_1120 => ce_1120_sg_x5,
      ce_2240 => ce_2240_sg_x5,
      ch_in => register1_q_net_x6,
      clk_1120 => clk_1120_sg_x5,
      clk_2240 => clk_2240_sg_x5,
      din => register4_q_net_x1,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_CORDIC"

entity fofb_cordic_entity_fad57e49ce is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ch_in: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(24 downto 0);
    q_in: in std_logic_vector(24 downto 0);
    valid_in: in std_logic;
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tddm_tbt_cordic0: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic0_x0: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic0_x1: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic0_x2: out std_logic_vector(23 downto 0)
  );
end fofb_cordic_entity_fad57e49ce;

architecture structural of fofb_cordic_entity_fad57e49ce is
  signal ce_1120_sg_x6: std_logic;
  signal ce_2240_sg_x6: std_logic;
  signal clk_1120_sg_x6: std_logic;
  signal clk_2240_sg_x6: std_logic;
  signal delay_q_net_x0: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tdata_phase_net: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tuser_cartesian_tuser_net: std_logic;
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register1_q_net_x7: std_logic;
  signal register4_q_net_x1: std_logic_vector(23 downto 0);
  signal register5_q_net_x5: std_logic_vector(23 downto 0);
  signal register_q_net_x1: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1120_sg_x6 <= ce_1120;
  ce_2240_sg_x6 <= ce_2240;
  delay_q_net_x0 <= ch_in;
  clk_1120_sg_x6 <= clk_1120;
  clk_2240_sg_x6 <= clk_2240;
  register_q_net_x2 <= i_in;
  register_q_net_x1 <= q_in;
  register1_q_net_x0 <= valid_in;
  amp_out <= register5_q_net_x5;
  ch_out <= register1_q_net_x7;
  tddm_tbt_cordic0 <= down_sample1_q_net_x4;
  tddm_tbt_cordic0_x0 <= down_sample2_q_net_x4;
  tddm_tbt_cordic0_x1 <= down_sample1_q_net_x5;
  tddm_tbt_cordic0_x2 <= down_sample2_q_net_x5;

  rect2pol: entity work.xlcordic_3fb964e2f71602f328fdd11ab57d7304
    port map (
      ce => ce_1120_sg_x6,
      clk => clk_1120_sg_x6,
      s_axis_cartesian_tdata_imag => register_q_net_x1,
      s_axis_cartesian_tdata_real => register_q_net_x2,
      s_axis_cartesian_tuser_user(0) => delay_q_net_x0,
      s_axis_cartesian_tvalid => register1_q_net_x0,
      m_axis_dout_tdata_phase => rect2pol_m_axis_dout_tdata_phase_net,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tuser_cartesian_tuser(0) => rect2pol_m_axis_dout_tuser_cartesian_tuser_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1120_sg_x6,
      clk => clk_1120_sg_x6,
      d(0) => rect2pol_m_axis_dout_tuser_cartesian_tuser_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q(0) => register1_q_net_x7
    );

  register4: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x6,
      clk => clk_1120_sg_x6,
      d => reinterpret2_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register4_q_net_x1
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x6,
      clk => clk_1120_sg_x6,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x5
    );

  reinterpret2: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_phase_net,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

  tddm_tbt_cordic0_38de3613fe: entity work.tddm_tbt_cordic0_entity_38de3613fe
    port map (
      ce_1120 => ce_1120_sg_x6,
      ce_2240 => ce_2240_sg_x6,
      clk_1120 => clk_1120_sg_x6,
      clk_2240 => clk_2240_sg_x6,
      fofb_cordic_ch_in => register1_q_net_x7,
      fofb_cordic_din => register5_q_net_x5,
      fofb_cordic_pin => register4_q_net_x1,
      fofb_cordic_data0_out => down_sample2_q_net_x4,
      fofb_cordic_data1_out => down_sample1_q_net_x4,
      fofb_cordic_phase0_out => down_sample2_q_net_x5,
      fofb_cordic_phase1_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp/Reg"

entity reg_entity_cf7aa296b2 is
  port (
    ce_1120: in std_logic;
    clk_1120: in std_logic;
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(23 downto 0)
  );
end reg_entity_cf7aa296b2;

architecture structural of reg_entity_cf7aa296b2 is
  signal ce_1120_sg_x7: std_logic;
  signal clk_1120_sg_x7: std_logic;
  signal convert_dout_net: std_logic_vector(23 downto 0);
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(24 downto 0);

begin
  ce_1120_sg_x7 <= ce_1120;
  clk_1120_sg_x7 <= clk_1120;
  register_q_net_x2 <= din;
  dout <= register_q_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 23,
      din_width => 25,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1120_sg_x7,
      clk => clk_1120_sg_x7,
      clr => '0',
      din => reinterpret2_output_port_net,
      en => "1",
      dout => convert_dout_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x7,
      clk => clk_1120_sg_x7,
      d => convert_dout_net,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

  reinterpret2: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => register_q_net_x2,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp/TDDM_fofb_cic0"

entity tddm_fofb_cic0_entity_6b909292ff is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    fofb_ch_in: in std_logic;
    fofb_i_in: in std_logic_vector(23 downto 0);
    fofb_q_in: in std_logic_vector(23 downto 0);
    cic_fofb_ch0_i_out: out std_logic_vector(23 downto 0);
    cic_fofb_ch0_q_out: out std_logic_vector(23 downto 0);
    cic_fofb_ch1_i_out: out std_logic_vector(23 downto 0);
    cic_fofb_ch1_q_out: out std_logic_vector(23 downto 0)
  );
end tddm_fofb_cic0_entity_6b909292ff;

architecture structural of tddm_fofb_cic0_entity_6b909292ff is
  signal ce_1120_sg_x11: std_logic;
  signal ce_2240_sg_x9: std_logic;
  signal clk_1120_sg_x11: std_logic;
  signal clk_2240_sg_x9: std_logic;
  signal delay_q_net_x3: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal register_q_net_x3: std_logic_vector(23 downto 0);
  signal register_q_net_x4: std_logic_vector(23 downto 0);

begin
  ce_1120_sg_x11 <= ce_1120;
  ce_2240_sg_x9 <= ce_2240;
  clk_1120_sg_x11 <= clk_1120;
  clk_2240_sg_x9 <= clk_2240;
  delay_q_net_x3 <= fofb_ch_in;
  register_q_net_x4 <= fofb_i_in;
  register_q_net_x3 <= fofb_q_in;
  cic_fofb_ch0_i_out <= down_sample2_q_net_x2;
  cic_fofb_ch0_q_out <= down_sample2_q_net_x3;
  cic_fofb_ch1_i_out <= down_sample1_q_net_x2;
  cic_fofb_ch1_q_out <= down_sample1_q_net_x3;

  tddm_fofb_cic0_i_06b84397ec: entity work.tddm_fofb_amp0_entity_fd74c6ad6e
    port map (
      ce_1120 => ce_1120_sg_x11,
      ce_2240 => ce_2240_sg_x9,
      ch_in => delay_q_net_x3,
      clk_1120 => clk_1120_sg_x11,
      clk_2240 => clk_2240_sg_x9,
      din => register_q_net_x4,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_fofb_cic0_q_a6a1d7c301: entity work.tddm_fofb_amp0_entity_fd74c6ad6e
    port map (
      ce_1120 => ce_1120_sg_x11,
      ce_2240 => ce_2240_sg_x9,
      ch_in => delay_q_net_x3,
      clk_1120 => clk_1120_sg_x11,
      clk_2240 => clk_2240_sg_x9,
      din => register_q_net_x3,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp/cic_fofb/Reg"

entity reg_entity_71dd029fba is
  port (
    ce_1120: in std_logic;
    clk_1120: in std_logic;
    din: in std_logic_vector(57 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(24 downto 0)
  );
end reg_entity_71dd029fba;

architecture structural of reg_entity_71dd029fba is
  signal ce_1120_sg_x12: std_logic;
  signal cic_fofb_q_m_axis_data_tdata_data_net_x0: std_logic_vector(57 downto 0);
  signal cic_fofb_q_m_axis_data_tvalid_net_x0: std_logic;
  signal clk_1120_sg_x12: std_logic;
  signal convert_dout_net: std_logic_vector(24 downto 0);
  signal register_q_net_x3: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(57 downto 0);

begin
  ce_1120_sg_x12 <= ce_1120;
  clk_1120_sg_x12 <= clk_1120;
  cic_fofb_q_m_axis_data_tdata_data_net_x0 <= din;
  cic_fofb_q_m_axis_data_tvalid_net_x0 <= en;
  dout <= register_q_net_x3;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 56,
      din_width => 58,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1120_sg_x12,
      clk => clk_1120_sg_x12,
      clr => '0',
      din => reinterpret2_output_port_net,
      en => "1",
      dout => convert_dout_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x12,
      clk => clk_1120_sg_x12,
      d => convert_dout_net,
      en(0) => cic_fofb_q_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x3
    );

  reinterpret2: entity work.reinterpret_fa01b5fd95
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_fofb_q_m_axis_data_tdata_data_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp/cic_fofb/Reg1"

entity reg1_entity_b079f30e3c is
  port (
    ce_1120: in std_logic;
    clk_1120: in std_logic;
    din: in std_logic_vector(57 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(24 downto 0);
    valid_out: out std_logic
  );
end reg1_entity_b079f30e3c;

architecture structural of reg1_entity_b079f30e3c is
  signal ce_1120_sg_x13: std_logic;
  signal cic_fofb_i_m_axis_data_tdata_data_net_x0: std_logic_vector(57 downto 0);
  signal cic_fofb_i_m_axis_data_tvalid_net_x0: std_logic;
  signal clk_1120_sg_x13: std_logic;
  signal convert_dout_net: std_logic_vector(24 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register_q_net_x4: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(57 downto 0);

begin
  ce_1120_sg_x13 <= ce_1120;
  clk_1120_sg_x13 <= clk_1120;
  cic_fofb_i_m_axis_data_tdata_data_net_x0 <= din;
  cic_fofb_i_m_axis_data_tvalid_net_x0 <= en;
  dout <= register_q_net_x4;
  valid_out <= register1_q_net_x1;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 56,
      din_width => 58,
      dout_arith => 2,
      dout_bin_pt => 23,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1120_sg_x13,
      clk => clk_1120_sg_x13,
      clr => '0',
      din => reinterpret2_output_port_net,
      en => "1",
      dout => convert_dout_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1120_sg_x13,
      clk => clk_1120_sg_x13,
      d(0) => cic_fofb_i_m_axis_data_tvalid_net_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x1
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x13,
      clk => clk_1120_sg_x13,
      d => convert_dout_net,
      en(0) => cic_fofb_i_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x4
    );

  reinterpret2: entity work.reinterpret_fa01b5fd95
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => cic_fofb_i_m_axis_data_tdata_data_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp/cic_fofb"

entity cic_fofb_entity_2ed6a6e00c is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    cic_fofb_q_x0: out std_logic;
    i_out: out std_logic_vector(24 downto 0);
    q_out: out std_logic_vector(24 downto 0);
    valid_out: out std_logic
  );
end cic_fofb_entity_2ed6a6e00c;

architecture structural of cic_fofb_entity_2ed6a6e00c is
  signal ce_1120_sg_x14: std_logic;
  signal ce_1_sg_x5: std_logic;
  signal ce_logic_1_sg_x5: std_logic;
  signal cic_fofb_i_m_axis_data_tdata_data_net_x0: std_logic_vector(57 downto 0);
  signal cic_fofb_i_m_axis_data_tuser_chan_out_net: std_logic;
  signal cic_fofb_i_m_axis_data_tvalid_net_x0: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x0: std_logic;
  signal cic_fofb_q_m_axis_data_tdata_data_net_x0: std_logic_vector(57 downto 0);
  signal cic_fofb_q_m_axis_data_tvalid_net_x0: std_logic;
  signal clk_1120_sg_x14: std_logic;
  signal clk_1_sg_x5: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal delay_q_net_x4: std_logic;
  signal register1_q_net_x2: std_logic;
  signal register3_q_net_x0: std_logic;
  signal register4_q_net_x0: std_logic_vector(23 downto 0);
  signal register5_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x5: std_logic_vector(24 downto 0);
  signal register_q_net_x6: std_logic_vector(24 downto 0);
  signal relational2_op_net: std_logic;

begin
  ce_1_sg_x5 <= ce_1;
  ce_1120_sg_x14 <= ce_1120;
  ce_logic_1_sg_x5 <= ce_logic_1;
  register3_q_net_x0 <= ch_in;
  clk_1_sg_x5 <= clk_1;
  clk_1120_sg_x14 <= clk_1120;
  register4_q_net_x0 <= i_in;
  register5_q_net_x0 <= q_in;
  ch_out <= delay_q_net_x4;
  cic_fofb_q_x0 <= cic_fofb_q_event_tlast_missing_net_x0;
  i_out <= register_q_net_x6;
  q_out <= register_q_net_x5;
  valid_out <= register1_q_net_x2;

  cic_fofb_i: entity work.xlcic_compiler_2d3b496704eca3daaae85383d488a908
    port map (
      ce => ce_1_sg_x5,
      ce_1120 => ce_1120_sg_x14,
      ce_logic_1 => ce_logic_1_sg_x5,
      clk => clk_1_sg_x5,
      clk_1120 => clk_1120_sg_x14,
      clk_logic_1 => clk_1_sg_x5,
      s_axis_data_tdata_data => register4_q_net_x0,
      s_axis_data_tlast => relational2_op_net,
      m_axis_data_tdata_data => cic_fofb_i_m_axis_data_tdata_data_net_x0,
      m_axis_data_tuser_chan_out(0) => cic_fofb_i_m_axis_data_tuser_chan_out_net,
      m_axis_data_tvalid => cic_fofb_i_m_axis_data_tvalid_net_x0
    );

  cic_fofb_q: entity work.xlcic_compiler_2d3b496704eca3daaae85383d488a908
    port map (
      ce => ce_1_sg_x5,
      ce_1120 => ce_1120_sg_x14,
      ce_logic_1 => ce_logic_1_sg_x5,
      clk => clk_1_sg_x5,
      clk_1120 => clk_1120_sg_x14,
      clk_logic_1 => clk_1_sg_x5,
      s_axis_data_tdata_data => register5_q_net_x0,
      s_axis_data_tlast => relational2_op_net,
      event_tlast_missing => cic_fofb_q_event_tlast_missing_net_x0,
      m_axis_data_tdata_data => cic_fofb_q_m_axis_data_tdata_data_net_x0,
      m_axis_data_tvalid => cic_fofb_q_m_axis_data_tvalid_net_x0
    );

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1120_sg_x14,
      clk => clk_1120_sg_x14,
      d(0) => cic_fofb_i_m_axis_data_tuser_chan_out_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x4
    );

  reg1_b079f30e3c: entity work.reg1_entity_b079f30e3c
    port map (
      ce_1120 => ce_1120_sg_x14,
      clk_1120 => clk_1120_sg_x14,
      din => cic_fofb_i_m_axis_data_tdata_data_net_x0,
      en => cic_fofb_i_m_axis_data_tvalid_net_x0,
      dout => register_q_net_x6,
      valid_out => register1_q_net_x2
    );

  reg_71dd029fba: entity work.reg_entity_71dd029fba
    port map (
      ce_1120 => ce_1120_sg_x14,
      clk_1120 => clk_1120_sg_x14,
      din => cic_fofb_q_m_axis_data_tdata_data_net_x0,
      en => cic_fofb_q_m_axis_data_tvalid_net_x0,
      dout => register_q_net_x5
    );

  relational2: entity work.relational_d29d27b7b3
    port map (
      a(0) => register3_q_net_x0,
      b => constant1_op_net,
      ce => ce_1_sg_x5,
      clk => clk_1_sg_x5,
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0/FOFB_amp"

entity fofb_amp_entity_078cdb1842 is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    cic_fofb: out std_logic;
    i_out: out std_logic_vector(24 downto 0);
    q_out: out std_logic_vector(24 downto 0);
    tddm_fofb_cic0: out std_logic_vector(23 downto 0);
    tddm_fofb_cic0_x0: out std_logic_vector(23 downto 0);
    tddm_fofb_cic0_x1: out std_logic_vector(23 downto 0);
    tddm_fofb_cic0_x2: out std_logic_vector(23 downto 0);
    valid_out: out std_logic
  );
end fofb_amp_entity_078cdb1842;

architecture structural of fofb_amp_entity_078cdb1842 is
  signal ce_1120_sg_x15: std_logic;
  signal ce_1_sg_x6: std_logic;
  signal ce_2240_sg_x10: std_logic;
  signal ce_logic_1_sg_x6: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x1: std_logic;
  signal clk_1120_sg_x15: std_logic;
  signal clk_1_sg_x6: std_logic;
  signal clk_2240_sg_x10: std_logic;
  signal delay_q_net_x5: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register3_q_net_x1: std_logic;
  signal register4_q_net_x1: std_logic_vector(23 downto 0);
  signal register5_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x3: std_logic_vector(23 downto 0);
  signal register_q_net_x4: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(24 downto 0);
  signal register_q_net_x8: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x6 <= ce_1;
  ce_1120_sg_x15 <= ce_1120;
  ce_2240_sg_x10 <= ce_2240;
  ce_logic_1_sg_x6 <= ce_logic_1;
  register3_q_net_x1 <= ch_in;
  clk_1_sg_x6 <= clk_1;
  clk_1120_sg_x15 <= clk_1120;
  clk_2240_sg_x10 <= clk_2240;
  register4_q_net_x1 <= i_in;
  register5_q_net_x1 <= q_in;
  ch_out <= delay_q_net_x5;
  cic_fofb <= cic_fofb_q_event_tlast_missing_net_x1;
  i_out <= register_q_net_x8;
  q_out <= register_q_net_x7;
  tddm_fofb_cic0 <= down_sample1_q_net_x4;
  tddm_fofb_cic0_x0 <= down_sample2_q_net_x4;
  tddm_fofb_cic0_x1 <= down_sample1_q_net_x5;
  tddm_fofb_cic0_x2 <= down_sample2_q_net_x5;
  valid_out <= register1_q_net_x3;

  cic_fofb_2ed6a6e00c: entity work.cic_fofb_entity_2ed6a6e00c
    port map (
      ce_1 => ce_1_sg_x6,
      ce_1120 => ce_1120_sg_x15,
      ce_logic_1 => ce_logic_1_sg_x6,
      ch_in => register3_q_net_x1,
      clk_1 => clk_1_sg_x6,
      clk_1120 => clk_1120_sg_x15,
      i_in => register4_q_net_x1,
      q_in => register5_q_net_x1,
      ch_out => delay_q_net_x5,
      cic_fofb_q_x0 => cic_fofb_q_event_tlast_missing_net_x1,
      i_out => register_q_net_x8,
      q_out => register_q_net_x7,
      valid_out => register1_q_net_x3
    );

  reg1_6375e37e24: entity work.reg_entity_cf7aa296b2
    port map (
      ce_1120 => ce_1120_sg_x15,
      clk_1120 => clk_1120_sg_x15,
      din => register_q_net_x8,
      dout => register_q_net_x4
    );

  reg_cf7aa296b2: entity work.reg_entity_cf7aa296b2
    port map (
      ce_1120 => ce_1120_sg_x15,
      clk_1120 => clk_1120_sg_x15,
      din => register_q_net_x7,
      dout => register_q_net_x3
    );

  tddm_fofb_cic0_6b909292ff: entity work.tddm_fofb_cic0_entity_6b909292ff
    port map (
      ce_1120 => ce_1120_sg_x15,
      ce_2240 => ce_2240_sg_x10,
      clk_1120 => clk_1120_sg_x15,
      clk_2240 => clk_2240_sg_x10,
      fofb_ch_in => delay_q_net_x5,
      fofb_i_in => register_q_net_x4,
      fofb_q_in => register_q_net_x3,
      cic_fofb_ch0_i_out => down_sample2_q_net_x4,
      cic_fofb_ch0_q_out => down_sample2_q_net_x5,
      cic_fofb_ch1_i_out => down_sample1_q_net_x4,
      cic_fofb_ch1_q_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp0"

entity fofb_amp0_entity_95b23bfc2c is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    fofb_amp: out std_logic_vector(23 downto 0);
    fofb_amp_x0: out std_logic_vector(23 downto 0);
    fofb_amp_x1: out std_logic_vector(23 downto 0);
    fofb_amp_x2: out std_logic_vector(23 downto 0);
    fofb_amp_x3: out std_logic;
    fofb_cordic: out std_logic_vector(23 downto 0);
    fofb_cordic_x0: out std_logic_vector(23 downto 0);
    fofb_cordic_x1: out std_logic_vector(23 downto 0);
    fofb_cordic_x2: out std_logic_vector(23 downto 0)
  );
end fofb_amp0_entity_95b23bfc2c;

architecture structural of fofb_amp0_entity_95b23bfc2c is
  signal ce_1120_sg_x16: std_logic;
  signal ce_1_sg_x7: std_logic;
  signal ce_2240_sg_x11: std_logic;
  signal ce_logic_1_sg_x7: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x2: std_logic;
  signal clk_1120_sg_x16: std_logic;
  signal clk_1_sg_x7: std_logic;
  signal clk_2240_sg_x11: std_logic;
  signal delay_q_net_x5: std_logic;
  signal down_sample1_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x9: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x9: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x8: std_logic;
  signal register3_q_net_x2: std_logic;
  signal register4_q_net_x2: std_logic_vector(23 downto 0);
  signal register5_q_net_x2: std_logic_vector(23 downto 0);
  signal register5_q_net_x6: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(24 downto 0);
  signal register_q_net_x8: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x7 <= ce_1;
  ce_1120_sg_x16 <= ce_1120;
  ce_2240_sg_x11 <= ce_2240;
  ce_logic_1_sg_x7 <= ce_logic_1;
  register3_q_net_x2 <= ch_in;
  clk_1_sg_x7 <= clk_1;
  clk_1120_sg_x16 <= clk_1120;
  clk_2240_sg_x11 <= clk_2240;
  register4_q_net_x2 <= i_in;
  register5_q_net_x2 <= q_in;
  amp_out <= register5_q_net_x6;
  ch_out <= register1_q_net_x8;
  fofb_amp <= down_sample1_q_net_x10;
  fofb_amp_x0 <= down_sample2_q_net_x10;
  fofb_amp_x1 <= down_sample1_q_net_x11;
  fofb_amp_x2 <= down_sample2_q_net_x11;
  fofb_amp_x3 <= cic_fofb_q_event_tlast_missing_net_x2;
  fofb_cordic <= down_sample1_q_net_x8;
  fofb_cordic_x0 <= down_sample2_q_net_x8;
  fofb_cordic_x1 <= down_sample1_q_net_x9;
  fofb_cordic_x2 <= down_sample2_q_net_x9;

  fofb_amp_078cdb1842: entity work.fofb_amp_entity_078cdb1842
    port map (
      ce_1 => ce_1_sg_x7,
      ce_1120 => ce_1120_sg_x16,
      ce_2240 => ce_2240_sg_x11,
      ce_logic_1 => ce_logic_1_sg_x7,
      ch_in => register3_q_net_x2,
      clk_1 => clk_1_sg_x7,
      clk_1120 => clk_1120_sg_x16,
      clk_2240 => clk_2240_sg_x11,
      i_in => register4_q_net_x2,
      q_in => register5_q_net_x2,
      ch_out => delay_q_net_x5,
      cic_fofb => cic_fofb_q_event_tlast_missing_net_x2,
      i_out => register_q_net_x8,
      q_out => register_q_net_x7,
      tddm_fofb_cic0 => down_sample1_q_net_x10,
      tddm_fofb_cic0_x0 => down_sample2_q_net_x10,
      tddm_fofb_cic0_x1 => down_sample1_q_net_x11,
      tddm_fofb_cic0_x2 => down_sample2_q_net_x11,
      valid_out => register1_q_net_x3
    );

  fofb_cordic_fad57e49ce: entity work.fofb_cordic_entity_fad57e49ce
    port map (
      ce_1120 => ce_1120_sg_x16,
      ce_2240 => ce_2240_sg_x11,
      ch_in => delay_q_net_x5,
      clk_1120 => clk_1120_sg_x16,
      clk_2240 => clk_2240_sg_x11,
      i_in => register_q_net_x8,
      q_in => register_q_net_x7,
      valid_in => register1_q_net_x3,
      amp_out => register5_q_net_x6,
      ch_out => register1_q_net_x8,
      tddm_tbt_cordic0 => down_sample1_q_net_x8,
      tddm_tbt_cordic0_x0 => down_sample2_q_net_x8,
      tddm_tbt_cordic0_x1 => down_sample1_q_net_x9,
      tddm_tbt_cordic0_x2 => down_sample2_q_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp1/FOFB_CORDIC"

entity fofb_cordic_entity_e4c0810ec7 is
  port (
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ch_in: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(24 downto 0);
    q_in: in std_logic_vector(24 downto 0);
    valid_in: in std_logic;
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tddm_fofb_cordic1: out std_logic_vector(23 downto 0);
    tddm_fofb_cordic1_x0: out std_logic_vector(23 downto 0);
    tddm_fofb_cordic1_x1: out std_logic_vector(23 downto 0);
    tddm_fofb_cordic1_x2: out std_logic_vector(23 downto 0)
  );
end fofb_cordic_entity_e4c0810ec7;

architecture structural of fofb_cordic_entity_e4c0810ec7 is
  signal ce_1120_sg_x20: std_logic;
  signal ce_2240_sg_x15: std_logic;
  signal clk_1120_sg_x20: std_logic;
  signal clk_2240_sg_x15: std_logic;
  signal delay_q_net_x0: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tdata_phase_net: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tdata_real_net: std_logic_vector(23 downto 0);
  signal rect2pol_m_axis_dout_tuser_cartesian_tuser_net: std_logic;
  signal rect2pol_m_axis_dout_tvalid_net: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register1_q_net_x8: std_logic;
  signal register4_q_net_x1: std_logic_vector(23 downto 0);
  signal register5_q_net_x6: std_logic_vector(23 downto 0);
  signal register_q_net_x1: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1120_sg_x20 <= ce_1120;
  ce_2240_sg_x15 <= ce_2240;
  delay_q_net_x0 <= ch_in;
  clk_1120_sg_x20 <= clk_1120;
  clk_2240_sg_x15 <= clk_2240;
  register_q_net_x2 <= i_in;
  register_q_net_x1 <= q_in;
  register1_q_net_x0 <= valid_in;
  amp_out <= register5_q_net_x6;
  ch_out <= register1_q_net_x8;
  tddm_fofb_cordic1 <= down_sample1_q_net_x4;
  tddm_fofb_cordic1_x0 <= down_sample2_q_net_x4;
  tddm_fofb_cordic1_x1 <= down_sample1_q_net_x5;
  tddm_fofb_cordic1_x2 <= down_sample2_q_net_x5;

  rect2pol: entity work.xlcordic_3fb964e2f71602f328fdd11ab57d7304
    port map (
      ce => ce_1120_sg_x20,
      clk => clk_1120_sg_x20,
      s_axis_cartesian_tdata_imag => register_q_net_x1,
      s_axis_cartesian_tdata_real => register_q_net_x2,
      s_axis_cartesian_tuser_user(0) => delay_q_net_x0,
      s_axis_cartesian_tvalid => register1_q_net_x0,
      m_axis_dout_tdata_phase => rect2pol_m_axis_dout_tdata_phase_net,
      m_axis_dout_tdata_real => rect2pol_m_axis_dout_tdata_real_net,
      m_axis_dout_tuser_cartesian_tuser(0) => rect2pol_m_axis_dout_tuser_cartesian_tuser_net,
      m_axis_dout_tvalid => rect2pol_m_axis_dout_tvalid_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1120_sg_x20,
      clk => clk_1120_sg_x20,
      d(0) => rect2pol_m_axis_dout_tuser_cartesian_tuser_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q(0) => register1_q_net_x8
    );

  register4: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x20,
      clk => clk_1120_sg_x20,
      d => reinterpret2_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register4_q_net_x1
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1120_sg_x20,
      clk => clk_1120_sg_x20,
      d => reinterpret3_output_port_net,
      en(0) => rect2pol_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x6
    );

  reinterpret2: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_phase_net,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => rect2pol_m_axis_dout_tdata_real_net,
      output_port => reinterpret3_output_port_net
    );

  tddm_fofb_cordic1_77b64089dc: entity work.tddm_tbt_cordic0_entity_38de3613fe
    port map (
      ce_1120 => ce_1120_sg_x20,
      ce_2240 => ce_2240_sg_x15,
      clk_1120 => clk_1120_sg_x20,
      clk_2240 => clk_2240_sg_x15,
      fofb_cordic_ch_in => register1_q_net_x8,
      fofb_cordic_din => register5_q_net_x6,
      fofb_cordic_pin => register4_q_net_x1,
      fofb_cordic_data0_out => down_sample2_q_net_x4,
      fofb_cordic_data1_out => down_sample1_q_net_x4,
      fofb_cordic_phase0_out => down_sample2_q_net_x5,
      fofb_cordic_phase1_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp1/FOFB_amp"

entity fofb_amp_entity_f70fcc8ed9 is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    cic_fofb: out std_logic;
    i_out: out std_logic_vector(24 downto 0);
    q_out: out std_logic_vector(24 downto 0);
    tddm_fofb_cic1: out std_logic_vector(23 downto 0);
    tddm_fofb_cic1_x0: out std_logic_vector(23 downto 0);
    tddm_fofb_cic1_x1: out std_logic_vector(23 downto 0);
    tddm_fofb_cic1_x2: out std_logic_vector(23 downto 0);
    valid_out: out std_logic
  );
end fofb_amp_entity_f70fcc8ed9;

architecture structural of fofb_amp_entity_f70fcc8ed9 is
  signal ce_1120_sg_x29: std_logic;
  signal ce_1_sg_x9: std_logic;
  signal ce_2240_sg_x19: std_logic;
  signal ce_logic_1_sg_x9: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x1: std_logic;
  signal clk_1120_sg_x29: std_logic;
  signal clk_1_sg_x9: std_logic;
  signal clk_2240_sg_x19: std_logic;
  signal delay_q_net_x5: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register3_q_net_x1: std_logic;
  signal register4_q_net_x1: std_logic_vector(23 downto 0);
  signal register5_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x3: std_logic_vector(23 downto 0);
  signal register_q_net_x4: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(24 downto 0);
  signal register_q_net_x8: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x9 <= ce_1;
  ce_1120_sg_x29 <= ce_1120;
  ce_2240_sg_x19 <= ce_2240;
  ce_logic_1_sg_x9 <= ce_logic_1;
  register3_q_net_x1 <= ch_in;
  clk_1_sg_x9 <= clk_1;
  clk_1120_sg_x29 <= clk_1120;
  clk_2240_sg_x19 <= clk_2240;
  register4_q_net_x1 <= i_in;
  register5_q_net_x1 <= q_in;
  ch_out <= delay_q_net_x5;
  cic_fofb <= cic_fofb_q_event_tlast_missing_net_x1;
  i_out <= register_q_net_x8;
  q_out <= register_q_net_x7;
  tddm_fofb_cic1 <= down_sample1_q_net_x4;
  tddm_fofb_cic1_x0 <= down_sample2_q_net_x4;
  tddm_fofb_cic1_x1 <= down_sample1_q_net_x5;
  tddm_fofb_cic1_x2 <= down_sample2_q_net_x5;
  valid_out <= register1_q_net_x3;

  cic_fofb_579902476d: entity work.cic_fofb_entity_2ed6a6e00c
    port map (
      ce_1 => ce_1_sg_x9,
      ce_1120 => ce_1120_sg_x29,
      ce_logic_1 => ce_logic_1_sg_x9,
      ch_in => register3_q_net_x1,
      clk_1 => clk_1_sg_x9,
      clk_1120 => clk_1120_sg_x29,
      i_in => register4_q_net_x1,
      q_in => register5_q_net_x1,
      ch_out => delay_q_net_x5,
      cic_fofb_q_x0 => cic_fofb_q_event_tlast_missing_net_x1,
      i_out => register_q_net_x8,
      q_out => register_q_net_x7,
      valid_out => register1_q_net_x3
    );

  reg1_a06a1c33b5: entity work.reg_entity_cf7aa296b2
    port map (
      ce_1120 => ce_1120_sg_x29,
      clk_1120 => clk_1120_sg_x29,
      din => register_q_net_x8,
      dout => register_q_net_x4
    );

  reg_b669a3b118: entity work.reg_entity_cf7aa296b2
    port map (
      ce_1120 => ce_1120_sg_x29,
      clk_1120 => clk_1120_sg_x29,
      din => register_q_net_x7,
      dout => register_q_net_x3
    );

  tddm_fofb_cic1_4a640315a5: entity work.tddm_fofb_cic0_entity_6b909292ff
    port map (
      ce_1120 => ce_1120_sg_x29,
      ce_2240 => ce_2240_sg_x19,
      clk_1120 => clk_1120_sg_x29,
      clk_2240 => clk_2240_sg_x19,
      fofb_ch_in => delay_q_net_x5,
      fofb_i_in => register_q_net_x4,
      fofb_q_in => register_q_net_x3,
      cic_fofb_ch0_i_out => down_sample2_q_net_x4,
      cic_fofb_ch0_q_out => down_sample2_q_net_x5,
      cic_fofb_ch1_i_out => down_sample1_q_net_x4,
      cic_fofb_ch1_q_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp/fofb_amp1"

entity fofb_amp1_entity_a049562dde is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    fofb_amp: out std_logic_vector(23 downto 0);
    fofb_amp_x0: out std_logic_vector(23 downto 0);
    fofb_amp_x1: out std_logic_vector(23 downto 0);
    fofb_amp_x2: out std_logic_vector(23 downto 0);
    fofb_amp_x3: out std_logic;
    fofb_cordic: out std_logic_vector(23 downto 0);
    fofb_cordic_x0: out std_logic_vector(23 downto 0);
    fofb_cordic_x1: out std_logic_vector(23 downto 0);
    fofb_cordic_x2: out std_logic_vector(23 downto 0)
  );
end fofb_amp1_entity_a049562dde;

architecture structural of fofb_amp1_entity_a049562dde is
  signal ce_1120_sg_x30: std_logic;
  signal ce_1_sg_x10: std_logic;
  signal ce_2240_sg_x20: std_logic;
  signal ce_logic_1_sg_x10: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x2: std_logic;
  signal clk_1120_sg_x30: std_logic;
  signal clk_1_sg_x10: std_logic;
  signal clk_2240_sg_x20: std_logic;
  signal delay_q_net_x5: std_logic;
  signal down_sample1_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x9: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x9: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x9: std_logic;
  signal register3_q_net_x2: std_logic;
  signal register4_q_net_x2: std_logic_vector(23 downto 0);
  signal register5_q_net_x2: std_logic_vector(23 downto 0);
  signal register5_q_net_x7: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(24 downto 0);
  signal register_q_net_x8: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x10 <= ce_1;
  ce_1120_sg_x30 <= ce_1120;
  ce_2240_sg_x20 <= ce_2240;
  ce_logic_1_sg_x10 <= ce_logic_1;
  register3_q_net_x2 <= ch_in;
  clk_1_sg_x10 <= clk_1;
  clk_1120_sg_x30 <= clk_1120;
  clk_2240_sg_x20 <= clk_2240;
  register4_q_net_x2 <= i_in;
  register5_q_net_x2 <= q_in;
  amp_out <= register5_q_net_x7;
  ch_out <= register1_q_net_x9;
  fofb_amp <= down_sample1_q_net_x10;
  fofb_amp_x0 <= down_sample2_q_net_x10;
  fofb_amp_x1 <= down_sample1_q_net_x11;
  fofb_amp_x2 <= down_sample2_q_net_x11;
  fofb_amp_x3 <= cic_fofb_q_event_tlast_missing_net_x2;
  fofb_cordic <= down_sample1_q_net_x8;
  fofb_cordic_x0 <= down_sample2_q_net_x8;
  fofb_cordic_x1 <= down_sample1_q_net_x9;
  fofb_cordic_x2 <= down_sample2_q_net_x9;

  fofb_amp_f70fcc8ed9: entity work.fofb_amp_entity_f70fcc8ed9
    port map (
      ce_1 => ce_1_sg_x10,
      ce_1120 => ce_1120_sg_x30,
      ce_2240 => ce_2240_sg_x20,
      ce_logic_1 => ce_logic_1_sg_x10,
      ch_in => register3_q_net_x2,
      clk_1 => clk_1_sg_x10,
      clk_1120 => clk_1120_sg_x30,
      clk_2240 => clk_2240_sg_x20,
      i_in => register4_q_net_x2,
      q_in => register5_q_net_x2,
      ch_out => delay_q_net_x5,
      cic_fofb => cic_fofb_q_event_tlast_missing_net_x2,
      i_out => register_q_net_x8,
      q_out => register_q_net_x7,
      tddm_fofb_cic1 => down_sample1_q_net_x10,
      tddm_fofb_cic1_x0 => down_sample2_q_net_x10,
      tddm_fofb_cic1_x1 => down_sample1_q_net_x11,
      tddm_fofb_cic1_x2 => down_sample2_q_net_x11,
      valid_out => register1_q_net_x3
    );

  fofb_cordic_e4c0810ec7: entity work.fofb_cordic_entity_e4c0810ec7
    port map (
      ce_1120 => ce_1120_sg_x30,
      ce_2240 => ce_2240_sg_x20,
      ch_in => delay_q_net_x5,
      clk_1120 => clk_1120_sg_x30,
      clk_2240 => clk_2240_sg_x20,
      i_in => register_q_net_x8,
      q_in => register_q_net_x7,
      valid_in => register1_q_net_x3,
      amp_out => register5_q_net_x7,
      ch_out => register1_q_net_x9,
      tddm_fofb_cordic1 => down_sample1_q_net_x8,
      tddm_fofb_cordic1_x0 => down_sample2_q_net_x8,
      tddm_fofb_cordic1_x1 => down_sample1_q_net_x9,
      tddm_fofb_cordic1_x2 => down_sample2_q_net_x9
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/FOFB_amp"

entity fofb_amp_entity_8b25d4b0b6 is
  port (
    ce_1: in std_logic;
    ce_1120: in std_logic;
    ce_2240: in std_logic;
    ce_logic_1: in std_logic;
    ch_in0: in std_logic;
    ch_in1: in std_logic;
    clk_1: in std_logic;
    clk_1120: in std_logic;
    clk_2240: in std_logic;
    i_in0: in std_logic_vector(23 downto 0);
    i_in1: in std_logic_vector(23 downto 0);
    q_in0: in std_logic_vector(23 downto 0);
    q_in1: in std_logic_vector(23 downto 0);
    amp_out0: out std_logic_vector(23 downto 0);
    amp_out1: out std_logic_vector(23 downto 0);
    amp_out2: out std_logic_vector(23 downto 0);
    amp_out3: out std_logic_vector(23 downto 0);
    fofb_amp0: out std_logic_vector(23 downto 0);
    fofb_amp0_x0: out std_logic_vector(23 downto 0);
    fofb_amp0_x1: out std_logic_vector(23 downto 0);
    fofb_amp0_x2: out std_logic_vector(23 downto 0);
    fofb_amp0_x3: out std_logic_vector(23 downto 0);
    fofb_amp0_x4: out std_logic_vector(23 downto 0);
    fofb_amp0_x5: out std_logic_vector(23 downto 0);
    fofb_amp0_x6: out std_logic_vector(23 downto 0);
    fofb_amp0_x7: out std_logic;
    fofb_amp1: out std_logic_vector(23 downto 0);
    fofb_amp1_x0: out std_logic_vector(23 downto 0);
    fofb_amp1_x1: out std_logic_vector(23 downto 0);
    fofb_amp1_x2: out std_logic_vector(23 downto 0);
    fofb_amp1_x3: out std_logic_vector(23 downto 0);
    fofb_amp1_x4: out std_logic_vector(23 downto 0);
    fofb_amp1_x5: out std_logic_vector(23 downto 0);
    fofb_amp1_x6: out std_logic_vector(23 downto 0);
    fofb_amp1_x7: out std_logic
  );
end fofb_amp_entity_8b25d4b0b6;

architecture structural of fofb_amp_entity_8b25d4b0b6 is
  signal ce_1120_sg_x31: std_logic;
  signal ce_1_sg_x11: std_logic;
  signal ce_2240_sg_x21: std_logic;
  signal ce_logic_1_sg_x11: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x4: std_logic;
  signal cic_fofb_q_event_tlast_missing_net_x5: std_logic;
  signal clk_1120_sg_x31: std_logic;
  signal clk_1_sg_x11: std_logic;
  signal clk_2240_sg_x21: std_logic;
  signal down_sample1_q_net_x16: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x17: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x19: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x22: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x23: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x24: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x25: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x16: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x17: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x19: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x22: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x23: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x24: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x25: std_logic_vector(23 downto 0);
  signal register1_q_net_x8: std_logic;
  signal register1_q_net_x9: std_logic;
  signal register3_q_net_x4: std_logic;
  signal register3_q_net_x5: std_logic;
  signal register4_q_net_x4: std_logic_vector(23 downto 0);
  signal register4_q_net_x5: std_logic_vector(23 downto 0);
  signal register5_q_net_x4: std_logic_vector(23 downto 0);
  signal register5_q_net_x6: std_logic_vector(23 downto 0);
  signal register5_q_net_x7: std_logic_vector(23 downto 0);
  signal register5_q_net_x8: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x11 <= ce_1;
  ce_1120_sg_x31 <= ce_1120;
  ce_2240_sg_x21 <= ce_2240;
  ce_logic_1_sg_x11 <= ce_logic_1;
  register3_q_net_x4 <= ch_in0;
  register3_q_net_x5 <= ch_in1;
  clk_1_sg_x11 <= clk_1;
  clk_1120_sg_x31 <= clk_1120;
  clk_2240_sg_x21 <= clk_2240;
  register4_q_net_x4 <= i_in0;
  register4_q_net_x5 <= i_in1;
  register5_q_net_x4 <= q_in0;
  register5_q_net_x8 <= q_in1;
  amp_out0 <= down_sample2_q_net_x16;
  amp_out1 <= down_sample1_q_net_x16;
  amp_out2 <= down_sample2_q_net_x17;
  amp_out3 <= down_sample1_q_net_x17;
  fofb_amp0 <= down_sample1_q_net_x18;
  fofb_amp0_x0 <= down_sample2_q_net_x18;
  fofb_amp0_x1 <= down_sample1_q_net_x19;
  fofb_amp0_x2 <= down_sample2_q_net_x19;
  fofb_amp0_x3 <= down_sample1_q_net_x20;
  fofb_amp0_x4 <= down_sample2_q_net_x20;
  fofb_amp0_x5 <= down_sample1_q_net_x21;
  fofb_amp0_x6 <= down_sample2_q_net_x21;
  fofb_amp0_x7 <= cic_fofb_q_event_tlast_missing_net_x4;
  fofb_amp1 <= down_sample1_q_net_x22;
  fofb_amp1_x0 <= down_sample2_q_net_x22;
  fofb_amp1_x1 <= down_sample1_q_net_x23;
  fofb_amp1_x2 <= down_sample2_q_net_x23;
  fofb_amp1_x3 <= down_sample1_q_net_x24;
  fofb_amp1_x4 <= down_sample2_q_net_x24;
  fofb_amp1_x5 <= down_sample1_q_net_x25;
  fofb_amp1_x6 <= down_sample2_q_net_x25;
  fofb_amp1_x7 <= cic_fofb_q_event_tlast_missing_net_x5;

  fofb_amp0_95b23bfc2c: entity work.fofb_amp0_entity_95b23bfc2c
    port map (
      ce_1 => ce_1_sg_x11,
      ce_1120 => ce_1120_sg_x31,
      ce_2240 => ce_2240_sg_x21,
      ce_logic_1 => ce_logic_1_sg_x11,
      ch_in => register3_q_net_x4,
      clk_1 => clk_1_sg_x11,
      clk_1120 => clk_1120_sg_x31,
      clk_2240 => clk_2240_sg_x21,
      i_in => register4_q_net_x4,
      q_in => register5_q_net_x4,
      amp_out => register5_q_net_x6,
      ch_out => register1_q_net_x8,
      fofb_amp => down_sample1_q_net_x20,
      fofb_amp_x0 => down_sample2_q_net_x20,
      fofb_amp_x1 => down_sample1_q_net_x21,
      fofb_amp_x2 => down_sample2_q_net_x21,
      fofb_amp_x3 => cic_fofb_q_event_tlast_missing_net_x4,
      fofb_cordic => down_sample1_q_net_x18,
      fofb_cordic_x0 => down_sample2_q_net_x18,
      fofb_cordic_x1 => down_sample1_q_net_x19,
      fofb_cordic_x2 => down_sample2_q_net_x19
    );

  fofb_amp1_a049562dde: entity work.fofb_amp1_entity_a049562dde
    port map (
      ce_1 => ce_1_sg_x11,
      ce_1120 => ce_1120_sg_x31,
      ce_2240 => ce_2240_sg_x21,
      ce_logic_1 => ce_logic_1_sg_x11,
      ch_in => register3_q_net_x5,
      clk_1 => clk_1_sg_x11,
      clk_1120 => clk_1120_sg_x31,
      clk_2240 => clk_2240_sg_x21,
      i_in => register4_q_net_x5,
      q_in => register5_q_net_x8,
      amp_out => register5_q_net_x7,
      ch_out => register1_q_net_x9,
      fofb_amp => down_sample1_q_net_x24,
      fofb_amp_x0 => down_sample2_q_net_x24,
      fofb_amp_x1 => down_sample1_q_net_x25,
      fofb_amp_x2 => down_sample2_q_net_x25,
      fofb_amp_x3 => cic_fofb_q_event_tlast_missing_net_x5,
      fofb_cordic => down_sample1_q_net_x22,
      fofb_cordic_x0 => down_sample2_q_net_x22,
      fofb_cordic_x1 => down_sample1_q_net_x23,
      fofb_cordic_x2 => down_sample2_q_net_x23
    );

  tddm_fofb_amp_4ch_2cc521a83f: entity work.tddm_fofb_amp_4ch_entity_2cc521a83f
    port map (
      amp_in0 => register5_q_net_x6,
      amp_in1 => register5_q_net_x7,
      ce_1120 => ce_1120_sg_x31,
      ce_2240 => ce_2240_sg_x21,
      ch_in0 => register1_q_net_x8,
      ch_in1 => register1_q_net_x9,
      clk_1120 => clk_1120_sg_x31,
      clk_2240 => clk_2240_sg_x21,
      amp_out0 => down_sample2_q_net_x16,
      amp_out1 => down_sample1_q_net_x16,
      amp_out2 => down_sample2_q_net_x17,
      amp_out3 => down_sample1_q_net_x17
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/K_fofb_mult3/Cast_truncate1"

entity cast_truncate1_entity_56731b7870 is
  port (
    in1: in std_logic_vector(49 downto 0);
    out1: out std_logic_vector(25 downto 0)
  );
end cast_truncate1_entity_56731b7870;

architecture structural of cast_truncate1_entity_56731b7870 is
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);
  signal slice_y_net: std_logic_vector(25 downto 0);

begin
  kx_tbt_p_net_x0 <= in1;
  out1 <= reinterpret_output_port_net_x0;

  reinterpret: entity work.reinterpret_9934b94a22
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_y_net,
      output_port => reinterpret_output_port_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 49,
      x_width => 50,
      y_width => 26
    )
    port map (
      x => kx_tbt_p_net_x0,
      y => slice_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/K_fofb_mult3"

entity k_fofb_mult3_entity_697accc8e2 is
  port (
    ce_2: in std_logic;
    ce_2240: in std_logic;
    clk_2: in std_logic;
    clk_2240: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end k_fofb_mult3_entity_697accc8e2;

architecture structural of k_fofb_mult3_entity_697accc8e2 is
  signal assert10_dout_net_x0: std_logic;
  signal assert5_dout_net_x0: std_logic_vector(24 downto 0);
  signal ce_2240_sg_x22: std_logic;
  signal ce_2_sg_x5: std_logic;
  signal clk_2240_sg_x22: std_logic;
  signal clk_2_sg_x5: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal kx_i_net_x0: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x5 <= ce_2;
  ce_2240_sg_x22 <= ce_2240;
  clk_2_sg_x5 <= clk_2;
  clk_2240_sg_x22 <= clk_2240;
  assert5_dout_net_x0 <= in1;
  kx_i_net_x0 <= in2;
  assert10_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_56731b7870: entity work.cast_truncate1_entity_56731b7870
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_2240_sg_x22,
      clk => clk_2240_sg_x22,
      d(0) => assert10_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 24,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 0,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 24,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert5_dout_net_x0,
      b => kx_i_net_x0,
      ce => ce_2_sg_x5,
      clk => clk_2_sg_x5,
      clr => '0',
      core_ce => ce_2_sg_x5,
      core_clk => clk_2_sg_x5,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x5,
      clk => clk_2_sg_x5,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/K_monit_1_mult"

entity k_monit_1_mult_entity_016885a3ac is
  port (
    ce_2: in std_logic;
    ce_224000000: in std_logic;
    clk_2: in std_logic;
    clk_224000000: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end k_monit_1_mult_entity_016885a3ac;

architecture structural of k_monit_1_mult_entity_016885a3ac is
  signal ce_224000000_sg_x0: std_logic;
  signal ce_2_sg_x8: std_logic;
  signal clk_224000000_sg_x0: std_logic;
  signal clk_2_sg_x8: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal kx_i_net_x2: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);
  signal ufix_to_bool_dout_net_x0: std_logic;

begin
  ce_2_sg_x8 <= ce_2;
  ce_224000000_sg_x0 <= ce_224000000;
  clk_2_sg_x8 <= clk_2;
  clk_224000000_sg_x0 <= clk_224000000;
  reinterpret3_output_port_net_x0 <= in1;
  kx_i_net_x2 <= in2;
  ufix_to_bool_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_fe5c8d5ea5: entity work.cast_truncate1_entity_56731b7870
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_224000000_sg_x0,
      clk => clk_224000000_sg_x0,
      d(0) => ufix_to_bool_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 24,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 0,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 24,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => reinterpret3_output_port_net_x0,
      b => kx_i_net_x2,
      ce => ce_2_sg_x8,
      clk => clk_2_sg_x8,
      clr => '0',
      core_ce => ce_2_sg_x8,
      core_clk => clk_2_sg_x8,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x8,
      clk => clk_2_sg_x8,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/K_monit_mult3"

entity k_monit_mult3_entity_8a778fb5f4 is
  port (
    ce_2: in std_logic;
    ce_22400000: in std_logic;
    clk_2: in std_logic;
    clk_22400000: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end k_monit_mult3_entity_8a778fb5f4;

architecture structural of k_monit_mult3_entity_8a778fb5f4 is
  signal assert11_dout_net_x0: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x0: std_logic;
  signal ce_22400000_sg_x0: std_logic;
  signal ce_2_sg_x11: std_logic;
  signal clk_22400000_sg_x0: std_logic;
  signal clk_2_sg_x11: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal kx_i_net_x4: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x11 <= ce_2;
  ce_22400000_sg_x0 <= ce_22400000;
  clk_2_sg_x11 <= clk_2;
  clk_22400000_sg_x0 <= clk_22400000;
  assert11_dout_net_x0 <= in1;
  kx_i_net_x4 <= in2;
  assert12_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_47fd83104e: entity work.cast_truncate1_entity_56731b7870
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_22400000_sg_x0,
      clk => clk_22400000_sg_x0,
      d(0) => assert12_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 24,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 0,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 24,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert11_dout_net_x0,
      b => kx_i_net_x4,
      ce => ce_2_sg_x11,
      clk => clk_2_sg_x11,
      clr => '0',
      core_ce => ce_2_sg_x11,
      core_clk => clk_2_sg_x11,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x11,
      clk => clk_2_sg_x11,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/K_tbt_mult"

entity k_tbt_mult_entity_b8fafff255 is
  port (
    ce_2: in std_logic;
    ce_70: in std_logic;
    clk_2: in std_logic;
    clk_70: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end k_tbt_mult_entity_b8fafff255;

architecture structural of k_tbt_mult_entity_b8fafff255 is
  signal assert10_dout_net_x0: std_logic;
  signal assert5_dout_net_x0: std_logic_vector(24 downto 0);
  signal ce_2_sg_x14: std_logic;
  signal ce_70_sg_x0: std_logic;
  signal clk_2_sg_x14: std_logic;
  signal clk_70_sg_x0: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal kx_i_net_x6: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x14 <= ce_2;
  ce_70_sg_x0 <= ce_70;
  clk_2_sg_x14 <= clk_2;
  clk_70_sg_x0 <= clk_70;
  assert5_dout_net_x0 <= in1;
  kx_i_net_x6 <= in2;
  assert10_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_4592ea30ee: entity work.cast_truncate1_entity_56731b7870
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_70_sg_x0,
      clk => clk_70_sg_x0,
      d(0) => assert10_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 24,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 0,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 24,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert5_dout_net_x0,
      b => kx_i_net_x6,
      ce => ce_2_sg_x14,
      clk => clk_2_sg_x14,
      clr => '0',
      core_ce => ce_2_sg_x14,
      core_clk => clk_2_sg_x14,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x14,
      clk => clk_2_sg_x14,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Ksum_fofb_mult4/Cast_truncate1"

entity cast_truncate1_entity_18a9b21a64 is
  port (
    in1: in std_logic_vector(49 downto 0);
    out1: out std_logic_vector(25 downto 0)
  );
end cast_truncate1_entity_18a9b21a64;

architecture structural of cast_truncate1_entity_18a9b21a64 is
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);
  signal slice_y_net: std_logic_vector(25 downto 0);

begin
  kx_tbt_p_net_x0 <= in1;
  out1 <= reinterpret_output_port_net_x0;

  reinterpret: entity work.reinterpret_9934b94a22
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_y_net,
      output_port => reinterpret_output_port_net_x0
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 49,
      x_width => 50,
      y_width => 26
    )
    port map (
      x => kx_tbt_p_net_x0,
      y => slice_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Ksum_fofb_mult4"

entity ksum_fofb_mult4_entity_ac3ed97096 is
  port (
    ce_2: in std_logic;
    ce_2240: in std_logic;
    clk_2: in std_logic;
    clk_2240: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end ksum_fofb_mult4_entity_ac3ed97096;

architecture structural of ksum_fofb_mult4_entity_ac3ed97096 is
  signal assert11_dout_net_x0: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x0: std_logic;
  signal ce_2240_sg_x25: std_logic;
  signal ce_2_sg_x17: std_logic;
  signal clk_2240_sg_x25: std_logic;
  signal clk_2_sg_x17: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal ksum_i_net_x0: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x17 <= ce_2;
  ce_2240_sg_x25 <= ce_2240;
  clk_2_sg_x17 <= clk_2;
  clk_2240_sg_x25 <= clk_2240;
  assert11_dout_net_x0 <= in1;
  ksum_i_net_x0 <= in2;
  assert12_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_18a9b21a64: entity work.cast_truncate1_entity_18a9b21a64
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_2240_sg_x25,
      clk => clk_2240_sg_x25,
      d(0) => assert12_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 21,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 44,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert11_dout_net_x0,
      b => ksum_i_net_x0,
      ce => ce_2_sg_x17,
      clk => clk_2_sg_x17,
      clr => '0',
      core_ce => ce_2_sg_x17,
      core_clk => clk_2_sg_x17,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x17,
      clk => clk_2_sg_x17,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Ksum_monit_1_mult1"

entity ksum_monit_1_mult1_entity_c66dc07078 is
  port (
    ce_2: in std_logic;
    ce_224000000: in std_logic;
    clk_2: in std_logic;
    clk_224000000: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end ksum_monit_1_mult1_entity_c66dc07078;

architecture structural of ksum_monit_1_mult1_entity_c66dc07078 is
  signal ce_224000000_sg_x3: std_logic;
  signal ce_2_sg_x18: std_logic;
  signal clk_224000000_sg_x3: std_logic;
  signal clk_2_sg_x18: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal ksum_i_net_x1: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret4_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);
  signal ufix_to_bool3_dout_net_x0: std_logic;

begin
  ce_2_sg_x18 <= ce_2;
  ce_224000000_sg_x3 <= ce_224000000;
  clk_2_sg_x18 <= clk_2;
  clk_224000000_sg_x3 <= clk_224000000;
  reinterpret4_output_port_net_x0 <= in1;
  ksum_i_net_x1 <= in2;
  ufix_to_bool3_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_92cc22397d: entity work.cast_truncate1_entity_18a9b21a64
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_224000000_sg_x3,
      clk => clk_224000000_sg_x3,
      d(0) => ufix_to_bool3_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 21,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 44,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => reinterpret4_output_port_net_x0,
      b => ksum_i_net_x1,
      ce => ce_2_sg_x18,
      clk => clk_2_sg_x18,
      clr => '0',
      core_ce => ce_2_sg_x18,
      core_clk => clk_2_sg_x18,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x18,
      clk => clk_2_sg_x18,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Ksum_monit_mult2"

entity ksum_monit_mult2_entity_31877b6d2b is
  port (
    ce_2: in std_logic;
    ce_22400000: in std_logic;
    clk_2: in std_logic;
    clk_22400000: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end ksum_monit_mult2_entity_31877b6d2b;

architecture structural of ksum_monit_mult2_entity_31877b6d2b is
  signal assert10_dout_net_x0: std_logic;
  signal assert5_dout_net_x0: std_logic_vector(24 downto 0);
  signal ce_22400000_sg_x3: std_logic;
  signal ce_2_sg_x19: std_logic;
  signal clk_22400000_sg_x3: std_logic;
  signal clk_2_sg_x19: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal ksum_i_net_x2: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x19 <= ce_2;
  ce_22400000_sg_x3 <= ce_22400000;
  clk_2_sg_x19 <= clk_2;
  clk_22400000_sg_x3 <= clk_22400000;
  assert5_dout_net_x0 <= in1;
  ksum_i_net_x2 <= in2;
  assert10_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_4c5b033963: entity work.cast_truncate1_entity_18a9b21a64
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_22400000_sg_x3,
      clk => clk_22400000_sg_x3,
      d(0) => assert10_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 21,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 44,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert5_dout_net_x0,
      b => ksum_i_net_x2,
      ce => ce_2_sg_x19,
      clk => clk_2_sg_x19,
      clr => '0',
      core_ce => ce_2_sg_x19,
      core_clk => clk_2_sg_x19,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x19,
      clk => clk_2_sg_x19,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Ksum_tbt_mult3"

entity ksum_tbt_mult3_entity_e0be30d675 is
  port (
    ce_2: in std_logic;
    ce_70: in std_logic;
    clk_2: in std_logic;
    clk_70: in std_logic;
    in1: in std_logic_vector(24 downto 0);
    in2: in std_logic_vector(24 downto 0);
    vld_in: in std_logic;
    out1: out std_logic_vector(25 downto 0);
    vld_out: out std_logic
  );
end ksum_tbt_mult3_entity_e0be30d675;

architecture structural of ksum_tbt_mult3_entity_e0be30d675 is
  signal assert11_dout_net_x0: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x0: std_logic;
  signal ce_2_sg_x20: std_logic;
  signal ce_70_sg_x3: std_logic;
  signal clk_2_sg_x20: std_logic;
  signal clk_70_sg_x3: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal ksum_i_net_x3: std_logic_vector(24 downto 0);
  signal kx_tbt_p_net_x0: std_logic_vector(49 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(25 downto 0);

begin
  ce_2_sg_x20 <= ce_2;
  ce_70_sg_x3 <= ce_70;
  clk_2_sg_x20 <= clk_2;
  clk_70_sg_x3 <= clk_70;
  assert11_dout_net_x0 <= in1;
  ksum_i_net_x3 <= in2;
  assert12_dout_net_x0 <= vld_in;
  out1 <= register_q_net_x0;
  vld_out <= delay1_q_net_x0;

  cast_truncate1_91bc0d396f: entity work.cast_truncate1_entity_18a9b21a64
    port map (
      in1 => kx_tbt_p_net_x0,
      out1 => reinterpret_output_port_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 9,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_70_sg_x3,
      clk => clk_70_sg_x3,
      d(0) => assert12_dout_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  kx_tbt: entity work.xlmult
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 21,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 23,
      b_width => 25,
      c_a_type => 0,
      c_a_width => 25,
      c_b_type => 0,
      c_b_width => 25,
      c_baat => 25,
      c_output_width => 50,
      c_type => 0,
      core_name0 => "mult_11_2_7786f9df1b07f80e",
      extra_registers => 0,
      multsign => 2,
      overflow => 1,
      p_arith => xlSigned,
      p_bin_pt => 44,
      p_width => 50,
      quantization => 1
    )
    port map (
      a => assert11_dout_net_x0,
      b => ksum_i_net_x3,
      ce => ce_2_sg_x20,
      clk => clk_2_sg_x20,
      clr => '0',
      core_ce => ce_2_sg_x20,
      core_clk => clk_2_sg_x20,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => kx_tbt_p_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x20,
      clk => clk_2_sg_x20,
      d => reinterpret_output_port_net_x0,
      en => "1",
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer/CMixer_0/DataReg_En"

entity datareg_en_entity_5c82ef2965 is
  port (
    ce_2: in std_logic;
    clk_2: in std_logic;
    din: in std_logic_vector(23 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(23 downto 0);
    valid: out std_logic
  );
end datareg_en_entity_5c82ef2965;

architecture structural of datareg_en_entity_5c82ef2965 is
  signal ce_2_sg_x21: std_logic;
  signal clk_2_sg_x21: std_logic;
  signal constant11_op_net_x0: std_logic;
  signal constant12_op_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);

begin
  ce_2_sg_x21 <= ce_2;
  clk_2_sg_x21 <= clk_2;
  constant12_op_net_x0 <= din;
  constant11_op_net_x0 <= en;
  dout <= register_q_net_x0;
  valid <= register1_q_net_x0;

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_2_sg_x21,
      clk => clk_2_sg_x21,
      d(0) => constant11_op_net_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x21,
      clk => clk_2_sg_x21,
      d => constant12_op_net_x0,
      en(0) => constant11_op_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer/CMixer_0/DataReg_En1"

entity datareg_en1_entity_8d533fde9e is
  port (
    ce_1: in std_logic;
    clk_1: in std_logic;
    din: in std_logic_vector(23 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(23 downto 0)
  );
end datareg_en1_entity_8d533fde9e;

architecture structural of datareg_en1_entity_8d533fde9e is
  signal ce_1_sg_x12: std_logic;
  signal clk_1_sg_x12: std_logic;
  signal constant11_op_net_x1: std_logic;
  signal register_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x2: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x12 <= ce_1;
  clk_1_sg_x12 <= clk_1;
  register_q_net_x1 <= din;
  constant11_op_net_x1 <= en;
  dout <= register_q_net_x2;

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x12,
      clk => clk_1_sg_x12,
      d => register_q_net_x1,
      en(0) => constant11_op_net_x1,
      rst => "0",
      q => register_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer/CMixer_0"

entity cmixer_0_entity_f630e8d7ec is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    dds_cosine: in std_logic_vector(23 downto 0);
    dds_msine: in std_logic_vector(23 downto 0);
    dds_valid: in std_logic;
    din_i: in std_logic_vector(23 downto 0);
    din_q: in std_logic_vector(23 downto 0);
    en: in std_logic;
    ch_out: out std_logic;
    i_out: out std_logic_vector(23 downto 0);
    q_out: out std_logic_vector(23 downto 0)
  );
end cmixer_0_entity_f630e8d7ec;

architecture structural of cmixer_0_entity_f630e8d7ec is
  signal a_i: std_logic_vector(23 downto 0);
  signal a_r: std_logic_vector(23 downto 0);
  signal b_i: std_logic_vector(23 downto 0);
  signal b_r: std_logic_vector(23 downto 0);
  signal ce_1_sg_x13: std_logic;
  signal ce_2_sg_x22: std_logic;
  signal clk_1_sg_x13: std_logic;
  signal clk_2_sg_x22: std_logic;
  signal complexmult_m_axis_dout_tdata_imag_net: std_logic_vector(23 downto 0);
  signal complexmult_m_axis_dout_tdata_real_net: std_logic_vector(23 downto 0);
  signal complexmult_m_axis_dout_tuser_net: std_logic;
  signal complexmult_m_axis_dout_tvalid_net: std_logic;
  signal constant11_op_net_x2: std_logic;
  signal constant12_op_net_x1: std_logic_vector(23 downto 0);
  signal constant15_op_net_x0: std_logic;
  signal convert1_dout_net: std_logic_vector(23 downto 0);
  signal convert2_dout_net: std_logic_vector(23 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register1_q_net_x1: std_logic;
  signal register3_q_net_x5: std_logic;
  signal register4_q_net_x5: std_logic_vector(23 downto 0);
  signal register5_q_net_x5: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x2: std_logic_vector(23 downto 0);
  signal register_q_net_x6: std_logic_vector(23 downto 0);
  signal register_q_net_x7: std_logic_vector(23 downto 0);
  signal register_q_net_x8: std_logic_vector(23 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x13 <= ce_1;
  ce_2_sg_x22 <= ce_2;
  register1_q_net_x1 <= ch_in;
  clk_1_sg_x13 <= clk_1;
  clk_2_sg_x22 <= clk_2;
  register_q_net_x6 <= dds_cosine;
  register_q_net_x7 <= dds_msine;
  constant15_op_net_x0 <= dds_valid;
  register_q_net_x8 <= din_i;
  constant12_op_net_x1 <= din_q;
  constant11_op_net_x2 <= en;
  ch_out <= register3_q_net_x5;
  i_out <= register4_q_net_x5;
  q_out <= register5_q_net_x5;

  complexmult: entity work.xlcomplex_multiplier_456da30af0f77a480cf80f52b29b4396
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      s_axis_a_tdata_imag => a_i,
      s_axis_a_tdata_real => a_r,
      s_axis_a_tvalid => constant15_op_net_x0,
      s_axis_b_tdata_imag => b_i,
      s_axis_b_tdata_real => b_r,
      s_axis_b_tuser(0) => register_q_net,
      s_axis_b_tvalid => register1_q_net_x0,
      m_axis_dout_tdata_imag => complexmult_m_axis_dout_tdata_imag_net,
      m_axis_dout_tdata_real => complexmult_m_axis_dout_tdata_real_net,
      m_axis_dout_tuser(0) => complexmult_m_axis_dout_tuser_net,
      m_axis_dout_tvalid => complexmult_m_axis_dout_tvalid_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 19,
      din_width => 24,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      clr => '0',
      din => reinterpret1_output_port_net,
      en => "1",
      dout => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 19,
      din_width => 24,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert2_dout_net
    );

  datareg_en1_8d533fde9e: entity work.datareg_en1_entity_8d533fde9e
    port map (
      ce_1 => ce_1_sg_x13,
      clk_1 => clk_1_sg_x13,
      din => register_q_net_x8,
      en => constant11_op_net_x2,
      dout => register_q_net_x2
    );

  datareg_en_5c82ef2965: entity work.datareg_en_entity_5c82ef2965
    port map (
      ce_2 => ce_2_sg_x22,
      clk_2 => clk_2_sg_x22,
      din => constant12_op_net_x1,
      en => constant11_op_net_x2,
      dout => register_q_net_x0,
      valid => register1_q_net_x0
    );

  delay: entity work.delay_961b43f67a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => register_q_net_x0,
      q => b_i
    );

  delay1: entity work.delay_961b43f67a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d => register_q_net_x2,
      q => b_r
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d => register_q_net_x6,
      en(0) => constant15_op_net_x0,
      rst => "0",
      q => a_r
    );

  register2: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d => register_q_net_x7,
      en(0) => constant15_op_net_x0,
      rst => "0",
      q => a_i
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d(0) => complexmult_m_axis_dout_tuser_net,
      en(0) => complexmult_m_axis_dout_tvalid_net,
      rst => "0",
      q(0) => register3_q_net_x5
    );

  register4: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d => convert1_dout_net,
      en(0) => complexmult_m_axis_dout_tvalid_net,
      rst => "0",
      q => register4_q_net_x5
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d => convert2_dout_net,
      en(0) => complexmult_m_axis_dout_tvalid_net,
      rst => "0",
      q => register5_q_net_x5
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d(0) => register1_q_net_x1,
      en(0) => constant11_op_net_x2,
      rst => "0",
      q(0) => register_q_net
    );

  reinterpret: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => complexmult_m_axis_dout_tdata_imag_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => complexmult_m_axis_dout_tdata_real_net,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer/TDDM_Mixer/TDDM_Mixer0_i"

entity tddm_mixer0_i_entity_f95b8f24ad is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_mixer0_i_entity_f95b8f24ad;

architecture structural of tddm_mixer0_i_entity_f95b8f24ad is
  signal ce_1_sg_x16: std_logic;
  signal ce_2_sg_x25: std_logic;
  signal clk_1_sg_x16: std_logic;
  signal clk_2_sg_x25: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register3_q_net_x6: std_logic;
  signal register4_q_net_x6: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_1_sg_x16 <= ce_1;
  ce_2_sg_x25 <= ce_2;
  register3_q_net_x6 <= ch_in;
  clk_1_sg_x16 <= clk_1;
  clk_2_sg_x25 <= clk_2;
  register4_q_net_x6 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_2_sg_x25,
      dest_clk => clk_2_sg_x25,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x16,
      src_clk => clk_1_sg_x16,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_2_sg_x25,
      dest_clk => clk_2_sg_x25,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x16,
      src_clk => clk_1_sg_x16,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      d => register4_q_net_x6,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      d => register4_q_net_x6,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => register3_q_net_x6,
      b(0) => constant_op_net,
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_d29d27b7b3
    port map (
      a(0) => register3_q_net_x6,
      b => constant1_op_net,
      ce => ce_1_sg_x16,
      clk => clk_1_sg_x16,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer/TDDM_Mixer"

entity tddm_mixer_entity_8537ade7b6 is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    mix0_ch_in: in std_logic;
    mix0_i_in: in std_logic_vector(23 downto 0);
    mix0_q_in: in std_logic_vector(23 downto 0);
    mix1_ch_in: in std_logic;
    mix1_i_in: in std_logic_vector(23 downto 0);
    mix1_q_in: in std_logic_vector(23 downto 0);
    mix_ch0_i_out: out std_logic_vector(23 downto 0);
    mix_ch0_q_out: out std_logic_vector(23 downto 0);
    mix_ch1_i_out: out std_logic_vector(23 downto 0);
    mix_ch1_q_out: out std_logic_vector(23 downto 0);
    mix_ch2_i_out: out std_logic_vector(23 downto 0);
    mix_ch2_q_out: out std_logic_vector(23 downto 0);
    mix_ch3_i_out: out std_logic_vector(23 downto 0);
    mix_ch3_q_out: out std_logic_vector(23 downto 0)
  );
end tddm_mixer_entity_8537ade7b6;

architecture structural of tddm_mixer_entity_8537ade7b6 is
  signal ce_1_sg_x20: std_logic;
  signal ce_2_sg_x29: std_logic;
  signal clk_1_sg_x20: std_logic;
  signal clk_2_sg_x29: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x6: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x7: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x6: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x7: std_logic_vector(23 downto 0);
  signal register3_q_net_x10: std_logic;
  signal register3_q_net_x9: std_logic;
  signal register4_q_net_x8: std_logic_vector(23 downto 0);
  signal register4_q_net_x9: std_logic_vector(23 downto 0);
  signal register5_q_net_x11: std_logic_vector(23 downto 0);
  signal register5_q_net_x7: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x20 <= ce_1;
  ce_2_sg_x29 <= ce_2;
  clk_1_sg_x20 <= clk_1;
  clk_2_sg_x29 <= clk_2;
  register3_q_net_x9 <= mix0_ch_in;
  register4_q_net_x8 <= mix0_i_in;
  register5_q_net_x7 <= mix0_q_in;
  register3_q_net_x10 <= mix1_ch_in;
  register4_q_net_x9 <= mix1_i_in;
  register5_q_net_x11 <= mix1_q_in;
  mix_ch0_i_out <= down_sample2_q_net_x4;
  mix_ch0_q_out <= down_sample2_q_net_x5;
  mix_ch1_i_out <= down_sample1_q_net_x4;
  mix_ch1_q_out <= down_sample1_q_net_x5;
  mix_ch2_i_out <= down_sample2_q_net_x6;
  mix_ch2_q_out <= down_sample2_q_net_x7;
  mix_ch3_i_out <= down_sample1_q_net_x6;
  mix_ch3_q_out <= down_sample1_q_net_x7;

  tddm_mixer0_i_f95b8f24ad: entity work.tddm_mixer0_i_entity_f95b8f24ad
    port map (
      ce_1 => ce_1_sg_x20,
      ce_2 => ce_2_sg_x29,
      ch_in => register3_q_net_x9,
      clk_1 => clk_1_sg_x20,
      clk_2 => clk_2_sg_x29,
      din => register4_q_net_x8,
      dout_ch0 => down_sample2_q_net_x4,
      dout_ch1 => down_sample1_q_net_x4
    );

  tddm_mixer0_q_2c5e18f496: entity work.tddm_mixer0_i_entity_f95b8f24ad
    port map (
      ce_1 => ce_1_sg_x20,
      ce_2 => ce_2_sg_x29,
      ch_in => register3_q_net_x9,
      clk_1 => clk_1_sg_x20,
      clk_2 => clk_2_sg_x29,
      din => register5_q_net_x7,
      dout_ch0 => down_sample2_q_net_x5,
      dout_ch1 => down_sample1_q_net_x5
    );

  tddm_mixer1_i_1afc4ccdba: entity work.tddm_mixer0_i_entity_f95b8f24ad
    port map (
      ce_1 => ce_1_sg_x20,
      ce_2 => ce_2_sg_x29,
      ch_in => register3_q_net_x10,
      clk_1 => clk_1_sg_x20,
      clk_2 => clk_2_sg_x29,
      din => register4_q_net_x9,
      dout_ch0 => down_sample2_q_net_x6,
      dout_ch1 => down_sample1_q_net_x6
    );

  tddm_mixer1_q_ee4acbed30: entity work.tddm_mixer0_i_entity_f95b8f24ad
    port map (
      ce_1 => ce_1_sg_x20,
      ce_2 => ce_2_sg_x29,
      ch_in => register3_q_net_x10,
      clk_1 => clk_1_sg_x20,
      clk_2 => clk_2_sg_x29,
      din => register5_q_net_x11,
      dout_ch0 => down_sample2_q_net_x7,
      dout_ch1 => down_sample1_q_net_x7
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Mixer"

entity mixer_entity_a1cd828545 is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ch_in0: in std_logic;
    ch_in1: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    dds_cosine_0: in std_logic_vector(23 downto 0);
    dds_cosine_1: in std_logic_vector(23 downto 0);
    dds_msine_0: in std_logic_vector(23 downto 0);
    dds_msine_1: in std_logic_vector(23 downto 0);
    dds_valid_0: in std_logic;
    dds_valid_1: in std_logic;
    din0: in std_logic_vector(23 downto 0);
    din1: in std_logic_vector(23 downto 0);
    ch_out0: out std_logic;
    ch_out1: out std_logic;
    i_out0: out std_logic_vector(23 downto 0);
    i_out1: out std_logic_vector(23 downto 0);
    q_out0: out std_logic_vector(23 downto 0);
    q_out1: out std_logic_vector(23 downto 0);
    tddm_mixer: out std_logic_vector(23 downto 0);
    tddm_mixer_x0: out std_logic_vector(23 downto 0);
    tddm_mixer_x1: out std_logic_vector(23 downto 0);
    tddm_mixer_x2: out std_logic_vector(23 downto 0);
    tddm_mixer_x3: out std_logic_vector(23 downto 0);
    tddm_mixer_x4: out std_logic_vector(23 downto 0);
    tddm_mixer_x5: out std_logic_vector(23 downto 0);
    tddm_mixer_x6: out std_logic_vector(23 downto 0)
  );
end mixer_entity_a1cd828545;

architecture structural of mixer_entity_a1cd828545 is
  signal ce_1_sg_x21: std_logic;
  signal ce_2_sg_x30: std_logic;
  signal clk_1_sg_x21: std_logic;
  signal clk_2_sg_x30: std_logic;
  signal constant11_op_net_x2: std_logic;
  signal constant12_op_net_x1: std_logic_vector(23 downto 0);
  signal constant15_op_net_x1: std_logic;
  signal constant1_op_net_x2: std_logic;
  signal constant2_op_net_x1: std_logic_vector(23 downto 0);
  signal constant3_op_net_x1: std_logic;
  signal down_sample1_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x9: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x9: std_logic_vector(23 downto 0);
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x4: std_logic;
  signal register3_q_net_x11: std_logic;
  signal register3_q_net_x12: std_logic;
  signal register4_q_net_x10: std_logic_vector(23 downto 0);
  signal register4_q_net_x11: std_logic_vector(23 downto 0);
  signal register5_q_net_x12: std_logic_vector(23 downto 0);
  signal register5_q_net_x8: std_logic_vector(23 downto 0);
  signal register_q_net_x12: std_logic_vector(23 downto 0);
  signal register_q_net_x13: std_logic_vector(23 downto 0);
  signal register_q_net_x14: std_logic_vector(23 downto 0);
  signal register_q_net_x15: std_logic_vector(23 downto 0);
  signal register_q_net_x16: std_logic_vector(23 downto 0);
  signal register_q_net_x17: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x21 <= ce_1;
  ce_2_sg_x30 <= ce_2;
  register1_q_net_x3 <= ch_in0;
  register1_q_net_x4 <= ch_in1;
  clk_1_sg_x21 <= clk_1;
  clk_2_sg_x30 <= clk_2;
  register_q_net_x12 <= dds_cosine_0;
  register_q_net_x14 <= dds_cosine_1;
  register_q_net_x13 <= dds_msine_0;
  register_q_net_x15 <= dds_msine_1;
  constant15_op_net_x1 <= dds_valid_0;
  constant3_op_net_x1 <= dds_valid_1;
  register_q_net_x16 <= din0;
  register_q_net_x17 <= din1;
  ch_out0 <= register3_q_net_x11;
  ch_out1 <= register3_q_net_x12;
  i_out0 <= register4_q_net_x10;
  i_out1 <= register4_q_net_x11;
  q_out0 <= register5_q_net_x8;
  q_out1 <= register5_q_net_x12;
  tddm_mixer <= down_sample1_q_net_x8;
  tddm_mixer_x0 <= down_sample2_q_net_x8;
  tddm_mixer_x1 <= down_sample1_q_net_x9;
  tddm_mixer_x2 <= down_sample2_q_net_x9;
  tddm_mixer_x3 <= down_sample1_q_net_x10;
  tddm_mixer_x4 <= down_sample2_q_net_x10;
  tddm_mixer_x5 <= down_sample1_q_net_x11;
  tddm_mixer_x6 <= down_sample2_q_net_x11;

  cmixer_0_f630e8d7ec: entity work.cmixer_0_entity_f630e8d7ec
    port map (
      ce_1 => ce_1_sg_x21,
      ce_2 => ce_2_sg_x30,
      ch_in => register1_q_net_x3,
      clk_1 => clk_1_sg_x21,
      clk_2 => clk_2_sg_x30,
      dds_cosine => register_q_net_x12,
      dds_msine => register_q_net_x13,
      dds_valid => constant15_op_net_x1,
      din_i => register_q_net_x16,
      din_q => constant12_op_net_x1,
      en => constant11_op_net_x2,
      ch_out => register3_q_net_x11,
      i_out => register4_q_net_x10,
      q_out => register5_q_net_x8
    );

  cmixer_1_61bfc18f90: entity work.cmixer_0_entity_f630e8d7ec
    port map (
      ce_1 => ce_1_sg_x21,
      ce_2 => ce_2_sg_x30,
      ch_in => register1_q_net_x4,
      clk_1 => clk_1_sg_x21,
      clk_2 => clk_2_sg_x30,
      dds_cosine => register_q_net_x14,
      dds_msine => register_q_net_x15,
      dds_valid => constant3_op_net_x1,
      din_i => register_q_net_x17,
      din_q => constant2_op_net_x1,
      en => constant1_op_net_x2,
      ch_out => register3_q_net_x12,
      i_out => register4_q_net_x11,
      q_out => register5_q_net_x12
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net_x2
    );

  constant11: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant11_op_net_x2
    );

  constant12: entity work.constant_f394f3309c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant12_op_net_x1
    );

  constant2: entity work.constant_f394f3309c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net_x1
    );

  tddm_mixer_8537ade7b6: entity work.tddm_mixer_entity_8537ade7b6
    port map (
      ce_1 => ce_1_sg_x21,
      ce_2 => ce_2_sg_x30,
      clk_1 => clk_1_sg_x21,
      clk_2 => clk_2_sg_x30,
      mix0_ch_in => register3_q_net_x11,
      mix0_i_in => register4_q_net_x10,
      mix0_q_in => register5_q_net_x8,
      mix1_ch_in => register3_q_net_x12,
      mix1_i_in => register4_q_net_x11,
      mix1_q_in => register5_q_net_x12,
      mix_ch0_i_out => down_sample2_q_net_x8,
      mix_ch0_q_out => down_sample2_q_net_x9,
      mix_ch1_i_out => down_sample1_q_net_x8,
      mix_ch1_q_out => down_sample1_q_net_x9,
      mix_ch2_i_out => down_sample2_q_net_x10,
      mix_ch2_q_out => down_sample2_q_net_x11,
      mix_ch3_i_out => down_sample1_q_net_x10,
      mix_ch3_q_out => down_sample1_q_net_x11
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/Cast2/format1"

entity format1_entity_4e0a69646b is
  port (
    ce_5600000: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(23 downto 0)
  );
end format1_entity_4e0a69646b;

architecture structural of format1_entity_4e0a69646b is
  signal ce_5600000_sg_x0: std_logic;
  signal clk_5600000_sg_x0: std_logic;
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal monit_pfir_m_axis_data_tdata_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(24 downto 0);

begin
  ce_5600000_sg_x0 <= ce_5600000;
  clk_5600000_sg_x0 <= clk_5600000;
  monit_pfir_m_axis_data_tdata_net_x0 <= din;
  dout <= convert_dout_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 21,
      din_width => 25,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_5600000_sg_x0,
      clk => clk_5600000_sg_x0,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  reinterpret: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => monit_pfir_m_axis_data_tdata_net_x0,
      output_port => reinterpret_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/Cast2"

entity cast2_entity_4b7421c7c9 is
  port (
    ce_5600000: in std_logic;
    clk_5600000: in std_logic;
    data_in: in std_logic_vector(24 downto 0);
    en: in std_logic;
    out_x0: out std_logic_vector(23 downto 0)
  );
end cast2_entity_4b7421c7c9;

architecture structural of cast2_entity_4b7421c7c9 is
  signal ce_5600000_sg_x1: std_logic;
  signal clk_5600000_sg_x1: std_logic;
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal monit_pfir_m_axis_data_tdata_net_x1: std_logic_vector(24 downto 0);
  signal monit_pfir_m_axis_data_tvalid_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);

begin
  ce_5600000_sg_x1 <= ce_5600000;
  clk_5600000_sg_x1 <= clk_5600000;
  monit_pfir_m_axis_data_tdata_net_x1 <= data_in;
  monit_pfir_m_axis_data_tvalid_net_x0 <= en;
  out_x0 <= register_q_net_x0;

  format1_4e0a69646b: entity work.format1_entity_4e0a69646b
    port map (
      ce_5600000 => ce_5600000_sg_x1,
      clk_5600000 => clk_5600000_sg_x1,
      din => monit_pfir_m_axis_data_tdata_net_x1,
      dout => convert_dout_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_5600000_sg_x1,
      clk => clk_5600000_sg_x1,
      d => convert_dout_net_x0,
      en(0) => monit_pfir_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/Cast4/format1"

entity format1_entity_3cf61b0d44 is
  port (
    ce_2800000: in std_logic;
    clk_2800000: in std_logic;
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(23 downto 0)
  );
end format1_entity_3cf61b0d44;

architecture structural of format1_entity_3cf61b0d44 is
  signal ce_2800000_sg_x0: std_logic;
  signal clk_2800000_sg_x0: std_logic;
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal monit_cfir_m_axis_data_tdata_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(24 downto 0);

begin
  ce_2800000_sg_x0 <= ce_2800000;
  clk_2800000_sg_x0 <= clk_2800000;
  monit_cfir_m_axis_data_tdata_net_x0 <= din;
  dout <= convert_dout_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 21,
      din_width => 25,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_2800000_sg_x0,
      clk => clk_2800000_sg_x0,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  reinterpret: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => monit_cfir_m_axis_data_tdata_net_x0,
      output_port => reinterpret_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/Cast4"

entity cast4_entity_4ed908d7fc is
  port (
    ce_2800000: in std_logic;
    clk_2800000: in std_logic;
    data_in: in std_logic_vector(24 downto 0);
    en: in std_logic;
    out_x0: out std_logic_vector(23 downto 0)
  );
end cast4_entity_4ed908d7fc;

architecture structural of cast4_entity_4ed908d7fc is
  signal ce_2800000_sg_x1: std_logic;
  signal clk_2800000_sg_x1: std_logic;
  signal convert_dout_net_x0: std_logic_vector(23 downto 0);
  signal monit_cfir_m_axis_data_tdata_net_x1: std_logic_vector(24 downto 0);
  signal monit_cfir_m_axis_data_tvalid_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);

begin
  ce_2800000_sg_x1 <= ce_2800000;
  clk_2800000_sg_x1 <= clk_2800000;
  monit_cfir_m_axis_data_tdata_net_x1 <= data_in;
  monit_cfir_m_axis_data_tvalid_net_x0 <= en;
  out_x0 <= register_q_net_x0;

  format1_3cf61b0d44: entity work.format1_entity_3cf61b0d44
    port map (
      ce_2800000 => ce_2800000_sg_x1,
      clk_2800000 => clk_2800000_sg_x1,
      din => monit_cfir_m_axis_data_tdata_net_x1,
      dout => convert_dout_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_2800000_sg_x1,
      clk => clk_2800000_sg_x1,
      d => convert_dout_net_x0,
      en(0) => monit_cfir_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/Reg1"

entity reg1_entity_8661a44192 is
  port (
    ce_1400000: in std_logic;
    clk_1400000: in std_logic;
    din: in std_logic_vector(60 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(23 downto 0)
  );
end reg1_entity_8661a44192;

architecture structural of reg1_entity_8661a44192 is
  signal ce_1400000_sg_x0: std_logic;
  signal clk_1400000_sg_x0: std_logic;
  signal convert_dout_net: std_logic_vector(23 downto 0);
  signal monit_cic_m_axis_data_tdata_data_net_x0: std_logic_vector(60 downto 0);
  signal monit_cic_m_axis_data_tvalid_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(60 downto 0);

begin
  ce_1400000_sg_x0 <= ce_1400000;
  clk_1400000_sg_x0 <= clk_1400000;
  monit_cic_m_axis_data_tdata_data_net_x0 <= din;
  monit_cic_m_axis_data_tvalid_net_x0 <= en;
  dout <= register_q_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 59,
      din_width => 61,
      dout_arith => 2,
      dout_bin_pt => 22,
      dout_width => 24,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_1400000_sg_x0,
      clk => clk_1400000_sg_x0,
      clr => '0',
      din => reinterpret2_output_port_net,
      en => "1",
      dout => convert_dout_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1400000_sg_x0,
      clk => clk_1400000_sg_x0,
      d => convert_dout_net,
      en(0) => monit_cic_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

  reinterpret2: entity work.reinterpret_c88e29aa6b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => monit_cic_m_axis_data_tdata_data_net_x0,
      output_port => reinterpret2_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/TDDM_monit_amp_c/TDDM_monit_amp_c_int"

entity tddm_monit_amp_c_int_entity_554a834349 is
  port (
    ce_22400000: in std_logic;
    ce_5600000: in std_logic;
    ch_in: in std_logic_vector(1 downto 0);
    clk_22400000: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0);
    dout_ch2: out std_logic_vector(23 downto 0);
    dout_ch3: out std_logic_vector(23 downto 0)
  );
end tddm_monit_amp_c_int_entity_554a834349;

architecture structural of tddm_monit_amp_c_int_entity_554a834349 is
  signal ce_22400000_sg_x4: std_logic;
  signal ce_5600000_sg_x2: std_logic;
  signal clk_22400000_sg_x4: std_logic;
  signal clk_5600000_sg_x2: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal delay2_q_net_x0: std_logic_vector(1 downto 0);
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register2_q_net: std_logic_vector(23 downto 0);
  signal register3_q_net: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal register_q_net_x1: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_22400000_sg_x4 <= ce_22400000;
  ce_5600000_sg_x2 <= ce_5600000;
  delay2_q_net_x0 <= ch_in;
  clk_22400000_sg_x4 <= clk_22400000;
  clk_5600000_sg_x2 <= clk_5600000;
  register_q_net_x1 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;
  dout_ch2 <= down_sample3_q_net_x0;
  dout_ch3 <= down_sample4_q_net_x0;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant3: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant_x0: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_22400000_sg_x4,
      dest_clk => clk_22400000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5600000_sg_x2,
      src_clk => clk_5600000_sg_x2,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_22400000_sg_x4,
      dest_clk => clk_22400000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5600000_sg_x2,
      src_clk => clk_5600000_sg_x2,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  down_sample3: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register2_q_net,
      dest_ce => ce_22400000_sg_x4,
      dest_clk => clk_22400000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5600000_sg_x2,
      src_clk => clk_5600000_sg_x2,
      src_clr => '0',
      q => down_sample3_q_net_x0
    );

  down_sample4: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register3_q_net,
      dest_ce => ce_22400000_sg_x4,
      dest_clk => clk_22400000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5600000_sg_x2,
      src_clk => clk_5600000_sg_x2,
      src_clr => '0',
      q => down_sample4_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      d => register_q_net_x1,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      d => register_q_net_x1,
      en(0) => relational2_op_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      d => register_q_net_x1,
      en(0) => relational3_op_net,
      rst => "0",
      q => register3_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      d => register_q_net_x1,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_367321bc0c
    port map (
      a => delay2_q_net_x0,
      b => constant_op_net,
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_367321bc0c
    port map (
      a => delay2_q_net_x0,
      b => constant1_op_net,
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_367321bc0c
    port map (
      a => delay2_q_net_x0,
      b => constant3_op_net,
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_367321bc0c
    port map (
      a => delay2_q_net_x0,
      b => constant4_op_net,
      ce => ce_5600000_sg_x2,
      clk => clk_5600000_sg_x2,
      clr => '0',
      op(0) => relational3_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c/TDDM_monit_amp_c"

entity tddm_monit_amp_c_entity_5b2613eff7 is
  port (
    ce_22400000: in std_logic;
    ce_5600000: in std_logic;
    clk_22400000: in std_logic;
    clk_5600000: in std_logic;
    monit_ch_in: in std_logic_vector(1 downto 0);
    monit_din: in std_logic_vector(23 downto 0);
    monit_ch0_out: out std_logic_vector(23 downto 0);
    monit_ch1_out: out std_logic_vector(23 downto 0);
    monit_ch2_out: out std_logic_vector(23 downto 0);
    monit_ch3_out: out std_logic_vector(23 downto 0)
  );
end tddm_monit_amp_c_entity_5b2613eff7;

architecture structural of tddm_monit_amp_c_entity_5b2613eff7 is
  signal ce_22400000_sg_x5: std_logic;
  signal ce_5600000_sg_x3: std_logic;
  signal clk_22400000_sg_x5: std_logic;
  signal clk_5600000_sg_x3: std_logic;
  signal delay2_q_net_x1: std_logic_vector(1 downto 0);
  signal down_sample1_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x2: std_logic_vector(23 downto 0);

begin
  ce_22400000_sg_x5 <= ce_22400000;
  ce_5600000_sg_x3 <= ce_5600000;
  clk_22400000_sg_x5 <= clk_22400000;
  clk_5600000_sg_x3 <= clk_5600000;
  delay2_q_net_x1 <= monit_ch_in;
  register_q_net_x2 <= monit_din;
  monit_ch0_out <= down_sample2_q_net_x1;
  monit_ch1_out <= down_sample1_q_net_x1;
  monit_ch2_out <= down_sample3_q_net_x1;
  monit_ch3_out <= down_sample4_q_net_x1;

  tddm_monit_amp_c_int_554a834349: entity work.tddm_monit_amp_c_int_entity_554a834349
    port map (
      ce_22400000 => ce_22400000_sg_x5,
      ce_5600000 => ce_5600000_sg_x3,
      ch_in => delay2_q_net_x1,
      clk_22400000 => clk_22400000_sg_x5,
      clk_5600000 => clk_5600000_sg_x3,
      din => register_q_net_x2,
      dout_ch0 => down_sample2_q_net_x1,
      dout_ch1 => down_sample1_q_net_x1,
      dout_ch2 => down_sample3_q_net_x1,
      dout_ch3 => down_sample4_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/Monit_amp_c"

entity monit_amp_c_entity_c83793ea71 is
  port (
    ce_1: in std_logic;
    ce_1400000: in std_logic;
    ce_22400000: in std_logic;
    ce_2800000: in std_logic;
    ce_560: in std_logic;
    ce_5600000: in std_logic;
    ce_logic_1400000: in std_logic;
    ce_logic_2800000: in std_logic;
    ce_logic_560: in std_logic;
    ch_in: in std_logic_vector(1 downto 0);
    clk_1: in std_logic;
    clk_1400000: in std_logic;
    clk_22400000: in std_logic;
    clk_2800000: in std_logic;
    clk_560: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(23 downto 0);
    amp_out: out std_logic_vector(23 downto 0);
    ch_out_x1: out std_logic_vector(1 downto 0);
    monit_cfir_x0: out std_logic;
    monit_cic_x0: out std_logic;
    monit_pfir_x0: out std_logic;
    tddm_monit_amp_c: out std_logic_vector(23 downto 0);
    tddm_monit_amp_c_x0: out std_logic_vector(23 downto 0);
    tddm_monit_amp_c_x1: out std_logic_vector(23 downto 0);
    tddm_monit_amp_c_x2: out std_logic_vector(23 downto 0)
  );
end monit_amp_c_entity_c83793ea71;

architecture structural of monit_amp_c_entity_c83793ea71 is
  signal ce_1400000_sg_x1: std_logic;
  signal ce_1_sg_x22: std_logic;
  signal ce_22400000_sg_x6: std_logic;
  signal ce_2800000_sg_x2: std_logic;
  signal ce_5600000_sg_x4: std_logic;
  signal ce_560_sg_x0: std_logic;
  signal ce_logic_1400000_sg_x0: std_logic;
  signal ce_logic_2800000_sg_x0: std_logic;
  signal ce_logic_560_sg_x0: std_logic;
  signal ch_out_x0: std_logic_vector(1 downto 0);
  signal clk_1400000_sg_x1: std_logic;
  signal clk_1_sg_x22: std_logic;
  signal clk_22400000_sg_x6: std_logic;
  signal clk_2800000_sg_x2: std_logic;
  signal clk_5600000_sg_x4: std_logic;
  signal clk_560_sg_x0: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal delay1_q_net: std_logic_vector(23 downto 0);
  signal delay2_q_net_x2: std_logic_vector(1 downto 0);
  signal delay3_q_net: std_logic_vector(23 downto 0);
  signal delay_q_net: std_logic_vector(1 downto 0);
  signal dout_x0: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x2: std_logic_vector(23 downto 0);
  signal monit_cfir_event_s_data_chanid_incorrect_net_x0: std_logic;
  signal monit_cfir_m_axis_data_tdata_net_x1: std_logic_vector(24 downto 0);
  signal monit_cfir_m_axis_data_tuser_chanid_net: std_logic_vector(1 downto 0);
  signal monit_cfir_m_axis_data_tvalid_net_x0: std_logic;
  signal monit_cic_event_tlast_unexpected_net_x0: std_logic;
  signal monit_cic_m_axis_data_tdata_data_net_x0: std_logic_vector(60 downto 0);
  signal monit_cic_m_axis_data_tuser_chan_out_net: std_logic_vector(1 downto 0);
  signal monit_cic_m_axis_data_tvalid_net_x0: std_logic;
  signal monit_pfir_event_s_data_chanid_incorrect_net_x0: std_logic;
  signal monit_pfir_m_axis_data_tdata_net_x1: std_logic_vector(24 downto 0);
  signal monit_pfir_m_axis_data_tuser_chanid_net: std_logic_vector(1 downto 0);
  signal monit_pfir_m_axis_data_tvalid_net_x0: std_logic;
  signal register3_q_net: std_logic_vector(1 downto 0);
  signal register_q_net_x0: std_logic_vector(23 downto 0);
  signal register_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x3: std_logic_vector(23 downto 0);
  signal relational2_op_net: std_logic;

begin
  ce_1_sg_x22 <= ce_1;
  ce_1400000_sg_x1 <= ce_1400000;
  ce_22400000_sg_x6 <= ce_22400000;
  ce_2800000_sg_x2 <= ce_2800000;
  ce_560_sg_x0 <= ce_560;
  ce_5600000_sg_x4 <= ce_5600000;
  ce_logic_1400000_sg_x0 <= ce_logic_1400000;
  ce_logic_2800000_sg_x0 <= ce_logic_2800000;
  ce_logic_560_sg_x0 <= ce_logic_560;
  ch_out_x0 <= ch_in;
  clk_1_sg_x22 <= clk_1;
  clk_1400000_sg_x1 <= clk_1400000;
  clk_22400000_sg_x6 <= clk_22400000;
  clk_2800000_sg_x2 <= clk_2800000;
  clk_560_sg_x0 <= clk_560;
  clk_5600000_sg_x4 <= clk_5600000;
  dout_x0 <= din;
  amp_out <= register_q_net_x3;
  ch_out_x1 <= delay2_q_net_x2;
  monit_cfir_x0 <= monit_cfir_event_s_data_chanid_incorrect_net_x0;
  monit_cic_x0 <= monit_cic_event_tlast_unexpected_net_x0;
  monit_pfir_x0 <= monit_pfir_event_s_data_chanid_incorrect_net_x0;
  tddm_monit_amp_c <= down_sample1_q_net_x2;
  tddm_monit_amp_c_x0 <= down_sample2_q_net_x2;
  tddm_monit_amp_c_x1 <= down_sample3_q_net_x2;
  tddm_monit_amp_c_x2 <= down_sample4_q_net_x2;

  cast2_4b7421c7c9: entity work.cast2_entity_4b7421c7c9
    port map (
      ce_5600000 => ce_5600000_sg_x4,
      clk_5600000 => clk_5600000_sg_x4,
      data_in => monit_pfir_m_axis_data_tdata_net_x1,
      en => monit_pfir_m_axis_data_tvalid_net_x0,
      out_x0 => register_q_net_x3
    );

  cast4_4ed908d7fc: entity work.cast4_entity_4ed908d7fc
    port map (
      ce_2800000 => ce_2800000_sg_x2,
      clk_2800000 => clk_2800000_sg_x2,
      data_in => monit_cfir_m_axis_data_tdata_net_x1,
      en => monit_cfir_m_axis_data_tvalid_net_x0,
      out_x0 => register_q_net_x0
    );

  constant1: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 3,
      reg_retiming => 0,
      reset => 0,
      width => 2
    )
    port map (
      ce => ce_1400000_sg_x1,
      clk => clk_1400000_sg_x1,
      d => monit_cic_m_axis_data_tuser_chan_out_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 3,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_560_sg_x0,
      clk => clk_560_sg_x0,
      d => dout_x0,
      en => '1',
      rst => '1',
      q => delay1_q_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 2
    )
    port map (
      ce => ce_5600000_sg_x4,
      clk => clk_5600000_sg_x4,
      d => monit_pfir_m_axis_data_tuser_chanid_net,
      en => '1',
      rst => '1',
      q => delay2_q_net_x2
    );

  delay3: entity work.xldelay
    generic map (
      latency => 2,
      reg_retiming => 0,
      reset => 0,
      width => 24
    )
    port map (
      ce => ce_1400000_sg_x1,
      clk => clk_1400000_sg_x1,
      d => register_q_net_x1,
      en => '1',
      rst => '1',
      q => delay3_q_net
    );

  monit_cfir: entity work.xlfir_compiler_2acadf5a08d72e0ee15ce4e1ac741dc6
    port map (
      ce => ce_1_sg_x22,
      ce_1400000 => ce_1400000_sg_x1,
      ce_2800000 => ce_2800000_sg_x2,
      ce_logic_1400000 => ce_logic_1400000_sg_x0,
      clk => clk_1_sg_x22,
      clk_1400000 => clk_1400000_sg_x1,
      clk_2800000 => clk_2800000_sg_x2,
      clk_logic_1400000 => clk_1400000_sg_x1,
      s_axis_data_tdata => delay3_q_net,
      s_axis_data_tuser_chanid => delay_q_net,
      src_ce => ce_1400000_sg_x1,
      src_clk => clk_1400000_sg_x1,
      event_s_data_chanid_incorrect => monit_cfir_event_s_data_chanid_incorrect_net_x0,
      m_axis_data_tdata => monit_cfir_m_axis_data_tdata_net_x1,
      m_axis_data_tuser_chanid => monit_cfir_m_axis_data_tuser_chanid_net,
      m_axis_data_tvalid => monit_cfir_m_axis_data_tvalid_net_x0
    );

  monit_cic: entity work.xlcic_compiler_6efc67831a277bdb0701519c5a976f20
    port map (
      ce => ce_1_sg_x22,
      ce_1400000 => ce_1400000_sg_x1,
      ce_560 => ce_560_sg_x0,
      ce_logic_560 => ce_logic_560_sg_x0,
      clk => clk_1_sg_x22,
      clk_1400000 => clk_1400000_sg_x1,
      clk_560 => clk_560_sg_x0,
      clk_logic_560 => clk_560_sg_x0,
      s_axis_data_tdata_data => delay1_q_net,
      s_axis_data_tlast => relational2_op_net,
      event_tlast_unexpected => monit_cic_event_tlast_unexpected_net_x0,
      m_axis_data_tdata_data => monit_cic_m_axis_data_tdata_data_net_x0,
      m_axis_data_tuser_chan_out => monit_cic_m_axis_data_tuser_chan_out_net,
      m_axis_data_tvalid => monit_cic_m_axis_data_tvalid_net_x0
    );

  monit_pfir: entity work.xlfir_compiler_1da691037bdf8c1b85b3b4502d6e9610
    port map (
      ce => ce_1_sg_x22,
      ce_2800000 => ce_2800000_sg_x2,
      ce_5600000 => ce_5600000_sg_x4,
      ce_logic_2800000 => ce_logic_2800000_sg_x0,
      clk => clk_1_sg_x22,
      clk_2800000 => clk_2800000_sg_x2,
      clk_5600000 => clk_5600000_sg_x4,
      clk_logic_2800000 => clk_2800000_sg_x2,
      s_axis_data_tdata => register_q_net_x0,
      s_axis_data_tuser_chanid => register3_q_net,
      src_ce => ce_2800000_sg_x2,
      src_clk => clk_2800000_sg_x2,
      event_s_data_chanid_incorrect => monit_pfir_event_s_data_chanid_incorrect_net_x0,
      m_axis_data_tdata => monit_pfir_m_axis_data_tdata_net_x1,
      m_axis_data_tuser_chanid => monit_pfir_m_axis_data_tuser_chanid_net,
      m_axis_data_tvalid => monit_pfir_m_axis_data_tvalid_net_x0
    );

  reg1_8661a44192: entity work.reg1_entity_8661a44192
    port map (
      ce_1400000 => ce_1400000_sg_x1,
      clk_1400000 => clk_1400000_sg_x1,
      din => monit_cic_m_axis_data_tdata_data_net_x0,
      en => monit_cic_m_axis_data_tvalid_net_x0,
      dout => register_q_net_x1
    );

  register3: entity work.xlregister
    generic map (
      d_width => 2,
      init_value => b"00"
    )
    port map (
      ce => ce_2800000_sg_x2,
      clk => clk_2800000_sg_x2,
      d => monit_cfir_m_axis_data_tuser_chanid_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  relational2: entity work.relational_83ca2c6a3c
    port map (
      a => ch_out_x0,
      b => constant1_op_net,
      ce => ce_560_sg_x0,
      clk => clk_560_sg_x0,
      clr => '0',
      op(0) => relational2_op_net
    );

  tddm_monit_amp_c_5b2613eff7: entity work.tddm_monit_amp_c_entity_5b2613eff7
    port map (
      ce_22400000 => ce_22400000_sg_x6,
      ce_5600000 => ce_5600000_sg_x4,
      clk_22400000 => clk_22400000_sg_x6,
      clk_5600000 => clk_5600000_sg_x4,
      monit_ch_in => delay2_q_net_x2,
      monit_din => register_q_net_x3,
      monit_ch0_out => down_sample2_q_net_x2,
      monit_ch1_out => down_sample1_q_net_x2,
      monit_ch2_out => down_sample3_q_net_x2,
      monit_ch3_out => down_sample4_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp/TDDM_monit_amp_out"

entity tddm_monit_amp_out_entity_521eb373cc is
  port (
    ce_22400000: in std_logic;
    ce_5600000: in std_logic;
    clk_22400000: in std_logic;
    clk_5600000: in std_logic;
    monit_amp_ch_in: in std_logic_vector(1 downto 0);
    monit_amp_din: in std_logic_vector(23 downto 0);
    monit_amp_data0_out: out std_logic_vector(23 downto 0);
    monit_amp_data1_out: out std_logic_vector(23 downto 0);
    monit_amp_data2_out: out std_logic_vector(23 downto 0);
    monit_amp_data3_out: out std_logic_vector(23 downto 0)
  );
end tddm_monit_amp_out_entity_521eb373cc;

architecture structural of tddm_monit_amp_out_entity_521eb373cc is
  signal ce_22400000_sg_x8: std_logic;
  signal ce_5600000_sg_x6: std_logic;
  signal clk_22400000_sg_x8: std_logic;
  signal clk_5600000_sg_x6: std_logic;
  signal delay2_q_net_x4: std_logic_vector(1 downto 0);
  signal down_sample1_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x1: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x1: std_logic_vector(23 downto 0);
  signal register_q_net_x5: std_logic_vector(23 downto 0);

begin
  ce_22400000_sg_x8 <= ce_22400000;
  ce_5600000_sg_x6 <= ce_5600000;
  clk_22400000_sg_x8 <= clk_22400000;
  clk_5600000_sg_x6 <= clk_5600000;
  delay2_q_net_x4 <= monit_amp_ch_in;
  register_q_net_x5 <= monit_amp_din;
  monit_amp_data0_out <= down_sample2_q_net_x1;
  monit_amp_data1_out <= down_sample1_q_net_x1;
  monit_amp_data2_out <= down_sample3_q_net_x1;
  monit_amp_data3_out <= down_sample4_q_net_x1;

  tddm_monit_amp_out_int_b60196c7a6: entity work.tddm_monit_amp_c_int_entity_554a834349
    port map (
      ce_22400000 => ce_22400000_sg_x8,
      ce_5600000 => ce_5600000_sg_x6,
      ch_in => delay2_q_net_x4,
      clk_22400000 => clk_22400000_sg_x8,
      clk_5600000 => clk_5600000_sg_x6,
      din => register_q_net_x5,
      dout_ch0 => down_sample2_q_net_x1,
      dout_ch1 => down_sample1_q_net_x1,
      dout_ch2 => down_sample3_q_net_x1,
      dout_ch3 => down_sample4_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/Monit_amp"

entity monit_amp_entity_44da74e268 is
  port (
    ce_1: in std_logic;
    ce_1400000: in std_logic;
    ce_22400000: in std_logic;
    ce_2800000: in std_logic;
    ce_560: in std_logic;
    ce_5600000: in std_logic;
    ce_logic_1400000: in std_logic;
    ce_logic_2800000: in std_logic;
    ce_logic_560: in std_logic;
    ch_in: in std_logic_vector(1 downto 0);
    clk_1: in std_logic;
    clk_1400000: in std_logic;
    clk_22400000: in std_logic;
    clk_2800000: in std_logic;
    clk_560: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(23 downto 0);
    amp_out0: out std_logic_vector(23 downto 0);
    amp_out1: out std_logic_vector(23 downto 0);
    amp_out2: out std_logic_vector(23 downto 0);
    amp_out3: out std_logic_vector(23 downto 0);
    monit_amp_c: out std_logic_vector(23 downto 0);
    monit_amp_c_x0: out std_logic_vector(23 downto 0);
    monit_amp_c_x1: out std_logic_vector(23 downto 0);
    monit_amp_c_x2: out std_logic_vector(23 downto 0);
    monit_amp_c_x3: out std_logic;
    monit_amp_c_x4: out std_logic;
    monit_amp_c_x5: out std_logic
  );
end monit_amp_entity_44da74e268;

architecture structural of monit_amp_entity_44da74e268 is
  signal ce_1400000_sg_x2: std_logic;
  signal ce_1_sg_x23: std_logic;
  signal ce_22400000_sg_x9: std_logic;
  signal ce_2800000_sg_x3: std_logic;
  signal ce_5600000_sg_x7: std_logic;
  signal ce_560_sg_x1: std_logic;
  signal ce_logic_1400000_sg_x1: std_logic;
  signal ce_logic_2800000_sg_x1: std_logic;
  signal ce_logic_560_sg_x1: std_logic;
  signal ch_out_x1: std_logic_vector(1 downto 0);
  signal clk_1400000_sg_x2: std_logic;
  signal clk_1_sg_x23: std_logic;
  signal clk_22400000_sg_x9: std_logic;
  signal clk_2800000_sg_x3: std_logic;
  signal clk_5600000_sg_x7: std_logic;
  signal clk_560_sg_x1: std_logic;
  signal delay2_q_net_x4: std_logic_vector(1 downto 0);
  signal dout_x1: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x4: std_logic_vector(23 downto 0);
  signal monit_cfir_event_s_data_chanid_incorrect_net_x1: std_logic;
  signal monit_cic_event_tlast_unexpected_net_x1: std_logic;
  signal monit_pfir_event_s_data_chanid_incorrect_net_x1: std_logic;
  signal register_q_net_x5: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x23 <= ce_1;
  ce_1400000_sg_x2 <= ce_1400000;
  ce_22400000_sg_x9 <= ce_22400000;
  ce_2800000_sg_x3 <= ce_2800000;
  ce_560_sg_x1 <= ce_560;
  ce_5600000_sg_x7 <= ce_5600000;
  ce_logic_1400000_sg_x1 <= ce_logic_1400000;
  ce_logic_2800000_sg_x1 <= ce_logic_2800000;
  ce_logic_560_sg_x1 <= ce_logic_560;
  ch_out_x1 <= ch_in;
  clk_1_sg_x23 <= clk_1;
  clk_1400000_sg_x2 <= clk_1400000;
  clk_22400000_sg_x9 <= clk_22400000;
  clk_2800000_sg_x3 <= clk_2800000;
  clk_560_sg_x1 <= clk_560;
  clk_5600000_sg_x7 <= clk_5600000;
  dout_x1 <= din;
  amp_out0 <= down_sample2_q_net_x4;
  amp_out1 <= down_sample1_q_net_x4;
  amp_out2 <= down_sample3_q_net_x4;
  amp_out3 <= down_sample4_q_net_x4;
  monit_amp_c <= down_sample1_q_net_x3;
  monit_amp_c_x0 <= down_sample2_q_net_x3;
  monit_amp_c_x1 <= down_sample3_q_net_x3;
  monit_amp_c_x2 <= down_sample4_q_net_x3;
  monit_amp_c_x3 <= monit_cfir_event_s_data_chanid_incorrect_net_x1;
  monit_amp_c_x4 <= monit_cic_event_tlast_unexpected_net_x1;
  monit_amp_c_x5 <= monit_pfir_event_s_data_chanid_incorrect_net_x1;

  monit_amp_c_c83793ea71: entity work.monit_amp_c_entity_c83793ea71
    port map (
      ce_1 => ce_1_sg_x23,
      ce_1400000 => ce_1400000_sg_x2,
      ce_22400000 => ce_22400000_sg_x9,
      ce_2800000 => ce_2800000_sg_x3,
      ce_560 => ce_560_sg_x1,
      ce_5600000 => ce_5600000_sg_x7,
      ce_logic_1400000 => ce_logic_1400000_sg_x1,
      ce_logic_2800000 => ce_logic_2800000_sg_x1,
      ce_logic_560 => ce_logic_560_sg_x1,
      ch_in => ch_out_x1,
      clk_1 => clk_1_sg_x23,
      clk_1400000 => clk_1400000_sg_x2,
      clk_22400000 => clk_22400000_sg_x9,
      clk_2800000 => clk_2800000_sg_x3,
      clk_560 => clk_560_sg_x1,
      clk_5600000 => clk_5600000_sg_x7,
      din => dout_x1,
      amp_out => register_q_net_x5,
      ch_out_x1 => delay2_q_net_x4,
      monit_cfir_x0 => monit_cfir_event_s_data_chanid_incorrect_net_x1,
      monit_cic_x0 => monit_cic_event_tlast_unexpected_net_x1,
      monit_pfir_x0 => monit_pfir_event_s_data_chanid_incorrect_net_x1,
      tddm_monit_amp_c => down_sample1_q_net_x3,
      tddm_monit_amp_c_x0 => down_sample2_q_net_x3,
      tddm_monit_amp_c_x1 => down_sample3_q_net_x3,
      tddm_monit_amp_c_x2 => down_sample4_q_net_x3
    );

  tddm_monit_amp_out_521eb373cc: entity work.tddm_monit_amp_out_entity_521eb373cc
    port map (
      ce_22400000 => ce_22400000_sg_x9,
      ce_5600000 => ce_5600000_sg_x7,
      clk_22400000 => clk_22400000_sg_x9,
      clk_5600000 => clk_5600000_sg_x7,
      monit_amp_ch_in => delay2_q_net_x4,
      monit_amp_din => register_q_net_x5,
      monit_amp_data0_out => down_sample2_q_net_x4,
      monit_amp_data1_out => down_sample1_q_net_x4,
      monit_amp_data2_out => down_sample3_q_net_x4,
      monit_amp_data3_out => down_sample4_q_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_CORDIC/TDDM_tbt_cordic/TDDM_tbt_cordic"

entity tddm_tbt_cordic_entity_5b94be40c5 is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic_entity_5b94be40c5;

architecture structural of tddm_tbt_cordic_entity_5b94be40c5 is
  signal ce_35_sg_x0: std_logic;
  signal ce_70_sg_x4: std_logic;
  signal clk_35_sg_x0: std_logic;
  signal clk_70_sg_x4: std_logic;
  signal constant1_op_net: std_logic;
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal p_amp_out_x0: std_logic_vector(23 downto 0);
  signal p_ch_out_x0: std_logic;
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_35_sg_x0 <= ce_35;
  ce_70_sg_x4 <= ce_70;
  p_ch_out_x0 <= ch_in;
  clk_35_sg_x0 <= clk_35;
  clk_70_sg_x4 <= clk_70;
  p_amp_out_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_70_sg_x4,
      dest_clk => clk_70_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x0,
      src_clk => clk_35_sg_x0,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_70_sg_x4,
      dest_clk => clk_70_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x0,
      src_clk => clk_35_sg_x0,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      d => p_amp_out_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      d => p_amp_out_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => p_ch_out_x0,
      b(0) => constant_op_net,
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_a892e1bf40
    port map (
      a(0) => p_ch_out_x0,
      b(0) => constant1_op_net,
      ce => ce_35_sg_x0,
      clk => clk_35_sg_x0,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_CORDIC/TDDM_tbt_cordic/TDDM_tbt_cordic1"

entity tddm_tbt_cordic1_entity_d3f44a687c is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic1_entity_d3f44a687c;

architecture structural of tddm_tbt_cordic1_entity_d3f44a687c is
  signal ce_35_sg_x1: std_logic;
  signal ce_70_sg_x5: std_logic;
  signal clk_35_sg_x1: std_logic;
  signal clk_70_sg_x5: std_logic;
  signal constant1_op_net: std_logic;
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal p_ch_out_x1: std_logic;
  signal p_phase_out_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register_q_net: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_35_sg_x1 <= ce_35;
  ce_70_sg_x5 <= ce_70;
  p_ch_out_x1 <= ch_in;
  clk_35_sg_x1 <= clk_35;
  clk_70_sg_x5 <= clk_70;
  p_phase_out_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_70_sg_x5,
      dest_clk => clk_70_sg_x5,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x1,
      src_clk => clk_35_sg_x1,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_70_sg_x5,
      dest_clk => clk_70_sg_x5,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x1,
      src_clk => clk_35_sg_x1,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      d => p_phase_out_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      d => p_phase_out_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => p_ch_out_x1,
      b(0) => constant_op_net,
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_a892e1bf40
    port map (
      a(0) => p_ch_out_x1,
      b(0) => constant1_op_net,
      ce => ce_35_sg_x1,
      clk => clk_35_sg_x1,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_CORDIC/TDDM_tbt_cordic"

entity tddm_tbt_cordic_entity_18d3979a26 is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    tbt_cordic_ch_in: in std_logic;
    tbt_cordic_din: in std_logic_vector(23 downto 0);
    tbt_cordic_pin: in std_logic_vector(23 downto 0);
    tbt_cordic_data0_out: out std_logic_vector(23 downto 0);
    tbt_cordic_data1_out: out std_logic_vector(23 downto 0);
    tbt_cordic_phase0_out: out std_logic_vector(23 downto 0);
    tbt_cordic_phase1_out: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic_entity_18d3979a26;

architecture structural of tddm_tbt_cordic_entity_18d3979a26 is
  signal ce_35_sg_x2: std_logic;
  signal ce_70_sg_x6: std_logic;
  signal clk_35_sg_x2: std_logic;
  signal clk_70_sg_x6: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal p_amp_out_x1: std_logic_vector(23 downto 0);
  signal p_ch_out_x2: std_logic;
  signal p_phase_out_x1: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x2 <= ce_35;
  ce_70_sg_x6 <= ce_70;
  clk_35_sg_x2 <= clk_35;
  clk_70_sg_x6 <= clk_70;
  p_ch_out_x2 <= tbt_cordic_ch_in;
  p_amp_out_x1 <= tbt_cordic_din;
  p_phase_out_x1 <= tbt_cordic_pin;
  tbt_cordic_data0_out <= down_sample2_q_net_x2;
  tbt_cordic_data1_out <= down_sample1_q_net_x2;
  tbt_cordic_phase0_out <= down_sample2_q_net_x3;
  tbt_cordic_phase1_out <= down_sample1_q_net_x3;

  tddm_tbt_cordic1_d3f44a687c: entity work.tddm_tbt_cordic1_entity_d3f44a687c
    port map (
      ce_35 => ce_35_sg_x2,
      ce_70 => ce_70_sg_x6,
      ch_in => p_ch_out_x2,
      clk_35 => clk_35_sg_x2,
      clk_70 => clk_70_sg_x6,
      din => p_phase_out_x1,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

  tddm_tbt_cordic_5b94be40c5: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x2,
      ce_70 => ce_70_sg_x6,
      ch_in => p_ch_out_x2,
      clk_35 => clk_35_sg_x2,
      clk_70 => clk_70_sg_x6,
      din => p_amp_out_x1,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_CORDIC"

entity tbt_cordic_entity_232cb2e43e is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(24 downto 0);
    q_in: in std_logic_vector(24 downto 0);
    valid_in: in std_logic;
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tddm_tbt_cordic: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x0: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x1: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x2: out std_logic_vector(23 downto 0)
  );
end tbt_cordic_entity_232cb2e43e;

architecture structural of tbt_cordic_entity_232cb2e43e is
  signal ce_35_sg_x3: std_logic;
  signal ce_70_sg_x7: std_logic;
  signal clk_35_sg_x3: std_logic;
  signal clk_70_sg_x7: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal p_amp_out_x2: std_logic_vector(23 downto 0);
  signal p_ch_out_x3: std_logic;
  signal p_phase_out_x1: std_logic_vector(23 downto 0);
  signal phase: std_logic_vector(23 downto 0);
  signal ready: std_logic;
  signal real_x0: std_logic;
  signal register1_q_net_x0: std_logic_vector(24 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register3_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal reinterpret2_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(23 downto 0);
  signal valid_out: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x3 <= ce_35;
  ce_70_sg_x7 <= ce_70;
  register2_q_net_x0 <= ch_in;
  clk_35_sg_x3 <= clk_35;
  clk_70_sg_x7 <= clk_70;
  register3_q_net_x0 <= i_in;
  register1_q_net_x0 <= q_in;
  register6_q_net_x0 <= valid_in;
  amp_out <= p_amp_out_x2;
  ch_out <= p_ch_out_x3;
  tddm_tbt_cordic <= down_sample1_q_net_x4;
  tddm_tbt_cordic_x0 <= down_sample2_q_net_x4;
  tddm_tbt_cordic_x1 <= down_sample1_q_net_x5;
  tddm_tbt_cordic_x2 <= down_sample2_q_net_x5;

  rect2pol: entity work.xlcordic_3fb964e2f71602f328fdd11ab57d7304
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      s_axis_cartesian_tdata_imag => register1_q_net_x0,
      s_axis_cartesian_tdata_real => register3_q_net_x0,
      s_axis_cartesian_tuser_user(0) => register2_q_net_x0,
      s_axis_cartesian_tvalid => register6_q_net_x0,
      m_axis_dout_tdata_phase => valid_out,
      m_axis_dout_tdata_real => phase,
      m_axis_dout_tuser_cartesian_tuser(0) => real_x0,
      m_axis_dout_tvalid => ready
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      d(0) => real_x0,
      en(0) => ready,
      rst => "0",
      q(0) => p_ch_out_x3
    );

  register4: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      d => reinterpret2_output_port_net,
      en(0) => ready,
      rst => "0",
      q => p_phase_out_x1
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x3,
      clk => clk_35_sg_x3,
      d => reinterpret3_output_port_net,
      en(0) => ready,
      rst => "0",
      q => p_amp_out_x2
    );

  reinterpret2: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => valid_out,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => phase,
      output_port => reinterpret3_output_port_net
    );

  tddm_tbt_cordic_18d3979a26: entity work.tddm_tbt_cordic_entity_18d3979a26
    port map (
      ce_35 => ce_35_sg_x3,
      ce_70 => ce_70_sg_x7,
      clk_35 => clk_35_sg_x3,
      clk_70 => clk_70_sg_x7,
      tbt_cordic_ch_in => p_ch_out_x3,
      tbt_cordic_din => p_amp_out_x2,
      tbt_cordic_pin => p_phase_out_x1,
      tbt_cordic_data0_out => down_sample2_q_net_x4,
      tbt_cordic_data1_out => down_sample1_q_net_x4,
      tbt_cordic_phase0_out => down_sample2_q_net_x5,
      tbt_cordic_phase1_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_poly_decim/TDDM_TBT/TDDM_tbt_poly_i"

entity tddm_tbt_poly_i_entity_469601736c is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    din: in std_logic_vector(23 downto 0);
    dout_ch0: out std_logic_vector(23 downto 0);
    dout_ch1: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_poly_i_entity_469601736c;

architecture structural of tddm_tbt_poly_i_entity_469601736c is
  signal ce_35_sg_x4: std_logic;
  signal ce_70_sg_x8: std_logic;
  signal clk_35_sg_x4: std_logic;
  signal clk_70_sg_x8: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant_op_net: std_logic;
  signal down_sample1_q_net_x0: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(23 downto 0);
  signal register1_q_net: std_logic_vector(23 downto 0);
  signal register2_q_net_x1: std_logic;
  signal register_q_net: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(23 downto 0);
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_35_sg_x4 <= ce_35;
  ce_70_sg_x8 <= ce_70;
  register2_q_net_x1 <= ch_in;
  clk_35_sg_x4 <= clk_35;
  clk_70_sg_x8 <= clk_70;
  reinterpret_output_port_net_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_70_sg_x8,
      dest_clk => clk_70_sg_x8,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x4,
      src_clk => clk_35_sg_x4,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 2,
      latency => 1,
      phase => 1,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => register_q_net,
      dest_ce => ce_70_sg_x8,
      dest_clk => clk_70_sg_x8,
      dest_clr => '0',
      en => "1",
      src_ce => ce_35_sg_x4,
      src_clk => clk_35_sg_x4,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x4,
      clk => clk_35_sg_x4,
      d => reinterpret_output_port_net_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x4,
      clk => clk_35_sg_x4,
      d => reinterpret_output_port_net_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity work.relational_a892e1bf40
    port map (
      a(0) => register2_q_net_x1,
      b(0) => constant_op_net,
      ce => ce_35_sg_x4,
      clk => clk_35_sg_x4,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_d29d27b7b3
    port map (
      a(0) => register2_q_net_x1,
      b => constant1_op_net,
      ce => ce_35_sg_x4,
      clk => clk_35_sg_x4,
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_poly_decim/TDDM_TBT"

entity tddm_tbt_entity_9ac9f65b0b is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    tbt_ch_in: in std_logic;
    tbt_i_in: in std_logic_vector(23 downto 0);
    tbt_q_in: in std_logic_vector(23 downto 0);
    poly35_ch0_i_out: out std_logic_vector(23 downto 0);
    poly35_ch0_q_out: out std_logic_vector(23 downto 0);
    poly35_ch1_i_out: out std_logic_vector(23 downto 0);
    poly35_ch1_q_out: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_entity_9ac9f65b0b;

architecture structural of tddm_tbt_entity_9ac9f65b0b is
  signal ce_35_sg_x6: std_logic;
  signal ce_70_sg_x10: std_logic;
  signal clk_35_sg_x6: std_logic;
  signal clk_70_sg_x10: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal register2_q_net_x3: std_logic;
  signal reinterpret_output_port_net_x2: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net_x3: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x6 <= ce_35;
  ce_70_sg_x10 <= ce_70;
  clk_35_sg_x6 <= clk_35;
  clk_70_sg_x10 <= clk_70;
  register2_q_net_x3 <= tbt_ch_in;
  reinterpret_output_port_net_x3 <= tbt_i_in;
  reinterpret_output_port_net_x2 <= tbt_q_in;
  poly35_ch0_i_out <= down_sample2_q_net_x2;
  poly35_ch0_q_out <= down_sample2_q_net_x3;
  poly35_ch1_i_out <= down_sample1_q_net_x2;
  poly35_ch1_q_out <= down_sample1_q_net_x3;

  tddm_tbt_poly_i_469601736c: entity work.tddm_tbt_poly_i_entity_469601736c
    port map (
      ce_35 => ce_35_sg_x6,
      ce_70 => ce_70_sg_x10,
      ch_in => register2_q_net_x3,
      clk_35 => clk_35_sg_x6,
      clk_70 => clk_70_sg_x10,
      din => reinterpret_output_port_net_x3,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_tbt_poly_q_8011b4e29e: entity work.tddm_tbt_poly_i_entity_469601736c
    port map (
      ce_35 => ce_35_sg_x6,
      ce_70 => ce_70_sg_x10,
      ch_in => register2_q_net_x3,
      clk_35 => clk_35_sg_x6,
      clk_70 => clk_70_sg_x10,
      din => reinterpret_output_port_net_x2,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_poly_decim/Trunc"

entity trunc_entity_e5eda8a5ac is
  port (
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(23 downto 0)
  );
end trunc_entity_e5eda8a5ac;

architecture structural of trunc_entity_e5eda8a5ac is
  signal register1_q_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x3: std_logic_vector(23 downto 0);
  signal slice_y_net: std_logic_vector(23 downto 0);

begin
  register1_q_net_x1 <= din;
  dout <= reinterpret_output_port_net_x3;

  reinterpret: entity work.reinterpret_4bf1ad328a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_y_net,
      output_port => reinterpret_output_port_net_x3
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 24,
      x_width => 25,
      y_width => 24
    )
    port map (
      x => register1_q_net_x1,
      y => slice_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0/TBT_poly_decim"

entity tbt_poly_decim_entity_4477ec06c2 is
  port (
    ce_1: in std_logic;
    ce_35: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    i_out: out std_logic_vector(24 downto 0);
    q_out: out std_logic_vector(24 downto 0);
    tbt_poly_x0: out std_logic;
    tddm_tbt: out std_logic_vector(23 downto 0);
    tddm_tbt_x0: out std_logic_vector(23 downto 0);
    tddm_tbt_x1: out std_logic_vector(23 downto 0);
    tddm_tbt_x2: out std_logic_vector(23 downto 0);
    valid_out: out std_logic
  );
end tbt_poly_decim_entity_4477ec06c2;

architecture structural of tbt_poly_decim_entity_4477ec06c2 is
  signal ce_1_sg_x24: std_logic;
  signal ce_35_sg_x7: std_logic;
  signal ce_70_sg_x11: std_logic;
  signal ce_logic_1_sg_x12: std_logic;
  signal clk_1_sg_x24: std_logic;
  signal clk_35_sg_x7: std_logic;
  signal clk_70_sg_x11: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal register1_q_net_x2: std_logic_vector(24 downto 0);
  signal register2_q_net_x4: std_logic;
  signal register3_q_net_x12: std_logic;
  signal register3_q_net_x2: std_logic_vector(24 downto 0);
  signal register4_q_net_x11: std_logic_vector(23 downto 0);
  signal register5_q_net_x9: std_logic_vector(23 downto 0);
  signal register6_q_net_x1: std_logic;
  signal reinterpret1_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x3: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net_x4: std_logic_vector(23 downto 0);
  signal tbt_poly_event_s_data_chanid_incorrect_net_x0: std_logic;
  signal tbt_poly_m_axis_data_tdata_path0_net: std_logic_vector(24 downto 0);
  signal tbt_poly_m_axis_data_tdata_path1_net: std_logic_vector(24 downto 0);
  signal tbt_poly_m_axis_data_tuser_chanid_net: std_logic;
  signal tbt_poly_m_axis_data_tvalid_net: std_logic;

begin
  ce_1_sg_x24 <= ce_1;
  ce_35_sg_x7 <= ce_35;
  ce_70_sg_x11 <= ce_70;
  ce_logic_1_sg_x12 <= ce_logic_1;
  register3_q_net_x12 <= ch_in;
  clk_1_sg_x24 <= clk_1;
  clk_35_sg_x7 <= clk_35;
  clk_70_sg_x11 <= clk_70;
  register4_q_net_x11 <= i_in;
  register5_q_net_x9 <= q_in;
  ch_out <= register2_q_net_x4;
  i_out <= register3_q_net_x2;
  q_out <= register1_q_net_x2;
  tbt_poly_x0 <= tbt_poly_event_s_data_chanid_incorrect_net_x0;
  tddm_tbt <= down_sample1_q_net_x4;
  tddm_tbt_x0 <= down_sample2_q_net_x4;
  tddm_tbt_x1 <= down_sample1_q_net_x5;
  tddm_tbt_x2 <= down_sample2_q_net_x5;
  valid_out <= register6_q_net_x1;

  register1: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d => reinterpret_output_port_net,
      en(0) => tbt_poly_m_axis_data_tvalid_net,
      rst => "0",
      q => register1_q_net_x2
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d(0) => tbt_poly_m_axis_data_tuser_chanid_net,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x4
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d => reinterpret1_output_port_net,
      en(0) => tbt_poly_m_axis_data_tvalid_net,
      rst => "0",
      q => register3_q_net_x2
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x7,
      clk => clk_35_sg_x7,
      d(0) => tbt_poly_m_axis_data_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x1
    );

  reinterpret: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => tbt_poly_m_axis_data_tdata_path1_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => tbt_poly_m_axis_data_tdata_path0_net,
      output_port => reinterpret1_output_port_net
    );

  tbt_poly: entity work.xlfir_compiler_f7093b59b74f3d511e09195b077ec73c
    port map (
      ce => ce_1_sg_x24,
      ce_35 => ce_35_sg_x7,
      ce_logic_1 => ce_logic_1_sg_x12,
      clk => clk_1_sg_x24,
      clk_35 => clk_35_sg_x7,
      clk_logic_1 => clk_1_sg_x24,
      s_axis_data_tdata_path0 => register4_q_net_x11,
      s_axis_data_tdata_path1 => register5_q_net_x9,
      s_axis_data_tuser_chanid(0) => register3_q_net_x12,
      src_ce => ce_1_sg_x24,
      src_clk => clk_1_sg_x24,
      event_s_data_chanid_incorrect => tbt_poly_event_s_data_chanid_incorrect_net_x0,
      m_axis_data_tdata_path0 => tbt_poly_m_axis_data_tdata_path0_net,
      m_axis_data_tdata_path1 => tbt_poly_m_axis_data_tdata_path1_net,
      m_axis_data_tuser_chanid(0) => tbt_poly_m_axis_data_tuser_chanid_net,
      m_axis_data_tvalid => tbt_poly_m_axis_data_tvalid_net
    );

  tddm_tbt_9ac9f65b0b: entity work.tddm_tbt_entity_9ac9f65b0b
    port map (
      ce_35 => ce_35_sg_x7,
      ce_70 => ce_70_sg_x11,
      clk_35 => clk_35_sg_x7,
      clk_70 => clk_70_sg_x11,
      tbt_ch_in => register2_q_net_x4,
      tbt_i_in => reinterpret_output_port_net_x4,
      tbt_q_in => reinterpret_output_port_net_x3,
      poly35_ch0_i_out => down_sample2_q_net_x4,
      poly35_ch0_q_out => down_sample2_q_net_x5,
      poly35_ch1_i_out => down_sample1_q_net_x4,
      poly35_ch1_q_out => down_sample1_q_net_x5
    );

  trunc1_841a61ebcc: entity work.trunc_entity_e5eda8a5ac
    port map (
      din => register3_q_net_x2,
      dout => reinterpret_output_port_net_x4
    );

  trunc_e5eda8a5ac: entity work.trunc_entity_e5eda8a5ac
    port map (
      din => register1_q_net_x2,
      dout => reinterpret_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp0"

entity tbt_amp0_entity_88b1c45f0e is
  port (
    ce_1: in std_logic;
    ce_35: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tbt_cordic: out std_logic_vector(23 downto 0);
    tbt_cordic_x0: out std_logic_vector(23 downto 0);
    tbt_cordic_x1: out std_logic_vector(23 downto 0);
    tbt_cordic_x2: out std_logic_vector(23 downto 0);
    tbt_poly_decim: out std_logic;
    tbt_poly_decim_x0: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x1: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x2: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x3: out std_logic_vector(23 downto 0)
  );
end tbt_amp0_entity_88b1c45f0e;

architecture structural of tbt_amp0_entity_88b1c45f0e is
  signal ce_1_sg_x25: std_logic;
  signal ce_35_sg_x8: std_logic;
  signal ce_70_sg_x12: std_logic;
  signal ce_logic_1_sg_x13: std_logic;
  signal clk_1_sg_x25: std_logic;
  signal clk_35_sg_x8: std_logic;
  signal clk_70_sg_x12: std_logic;
  signal down_sample1_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x9: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x9: std_logic_vector(23 downto 0);
  signal p_amp_out_x3: std_logic_vector(23 downto 0);
  signal p_ch_out_x4: std_logic;
  signal register1_q_net_x2: std_logic_vector(24 downto 0);
  signal register2_q_net_x4: std_logic;
  signal register3_q_net_x13: std_logic;
  signal register3_q_net_x2: std_logic_vector(24 downto 0);
  signal register4_q_net_x12: std_logic_vector(23 downto 0);
  signal register5_q_net_x10: std_logic_vector(23 downto 0);
  signal register6_q_net_x1: std_logic;
  signal tbt_poly_event_s_data_chanid_incorrect_net_x1: std_logic;

begin
  ce_1_sg_x25 <= ce_1;
  ce_35_sg_x8 <= ce_35;
  ce_70_sg_x12 <= ce_70;
  ce_logic_1_sg_x13 <= ce_logic_1;
  register3_q_net_x13 <= ch_in;
  clk_1_sg_x25 <= clk_1;
  clk_35_sg_x8 <= clk_35;
  clk_70_sg_x12 <= clk_70;
  register4_q_net_x12 <= i_in;
  register5_q_net_x10 <= q_in;
  amp_out <= p_amp_out_x3;
  ch_out <= p_ch_out_x4;
  tbt_cordic <= down_sample1_q_net_x8;
  tbt_cordic_x0 <= down_sample2_q_net_x8;
  tbt_cordic_x1 <= down_sample1_q_net_x9;
  tbt_cordic_x2 <= down_sample2_q_net_x9;
  tbt_poly_decim <= tbt_poly_event_s_data_chanid_incorrect_net_x1;
  tbt_poly_decim_x0 <= down_sample1_q_net_x10;
  tbt_poly_decim_x1 <= down_sample2_q_net_x10;
  tbt_poly_decim_x2 <= down_sample1_q_net_x11;
  tbt_poly_decim_x3 <= down_sample2_q_net_x11;

  tbt_cordic_232cb2e43e: entity work.tbt_cordic_entity_232cb2e43e
    port map (
      ce_35 => ce_35_sg_x8,
      ce_70 => ce_70_sg_x12,
      ch_in => register2_q_net_x4,
      clk_35 => clk_35_sg_x8,
      clk_70 => clk_70_sg_x12,
      i_in => register3_q_net_x2,
      q_in => register1_q_net_x2,
      valid_in => register6_q_net_x1,
      amp_out => p_amp_out_x3,
      ch_out => p_ch_out_x4,
      tddm_tbt_cordic => down_sample1_q_net_x8,
      tddm_tbt_cordic_x0 => down_sample2_q_net_x8,
      tddm_tbt_cordic_x1 => down_sample1_q_net_x9,
      tddm_tbt_cordic_x2 => down_sample2_q_net_x9
    );

  tbt_poly_decim_4477ec06c2: entity work.tbt_poly_decim_entity_4477ec06c2
    port map (
      ce_1 => ce_1_sg_x25,
      ce_35 => ce_35_sg_x8,
      ce_70 => ce_70_sg_x12,
      ce_logic_1 => ce_logic_1_sg_x13,
      ch_in => register3_q_net_x13,
      clk_1 => clk_1_sg_x25,
      clk_35 => clk_35_sg_x8,
      clk_70 => clk_70_sg_x12,
      i_in => register4_q_net_x12,
      q_in => register5_q_net_x10,
      ch_out => register2_q_net_x4,
      i_out => register3_q_net_x2,
      q_out => register1_q_net_x2,
      tbt_poly_x0 => tbt_poly_event_s_data_chanid_incorrect_net_x1,
      tddm_tbt => down_sample1_q_net_x10,
      tddm_tbt_x0 => down_sample2_q_net_x10,
      tddm_tbt_x1 => down_sample1_q_net_x11,
      tddm_tbt_x2 => down_sample2_q_net_x11,
      valid_out => register6_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp1/TBT_CORDIC/TDDM_tbt_cordic"

entity tddm_tbt_cordic_entity_9e99bd206d is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    tbt_cordic_ch_in: in std_logic;
    tbt_cordic_din: in std_logic_vector(23 downto 0);
    tbt_cordic_pin: in std_logic_vector(23 downto 0);
    tbt_cordic_ch2_out: out std_logic_vector(23 downto 0);
    tbt_cordic_ch3_out: out std_logic_vector(23 downto 0);
    tbt_cordic_phase0_out: out std_logic_vector(23 downto 0);
    tbt_cordic_phase1_out: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_cordic_entity_9e99bd206d;

architecture structural of tddm_tbt_cordic_entity_9e99bd206d is
  signal ce_35_sg_x11: std_logic;
  signal ce_70_sg_x15: std_logic;
  signal clk_35_sg_x11: std_logic;
  signal clk_70_sg_x15: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal p_amp_out_x1: std_logic_vector(23 downto 0);
  signal p_ch_out_x2: std_logic;
  signal p_phase_out_x1: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x11 <= ce_35;
  ce_70_sg_x15 <= ce_70;
  clk_35_sg_x11 <= clk_35;
  clk_70_sg_x15 <= clk_70;
  p_ch_out_x2 <= tbt_cordic_ch_in;
  p_amp_out_x1 <= tbt_cordic_din;
  p_phase_out_x1 <= tbt_cordic_pin;
  tbt_cordic_ch2_out <= down_sample2_q_net_x2;
  tbt_cordic_ch3_out <= down_sample1_q_net_x2;
  tbt_cordic_phase0_out <= down_sample2_q_net_x3;
  tbt_cordic_phase1_out <= down_sample1_q_net_x3;

  tddm_tbt_cordic1_d22fbdac88: entity work.tddm_tbt_cordic1_entity_d3f44a687c
    port map (
      ce_35 => ce_35_sg_x11,
      ce_70 => ce_70_sg_x15,
      ch_in => p_ch_out_x2,
      clk_35 => clk_35_sg_x11,
      clk_70 => clk_70_sg_x15,
      din => p_phase_out_x1,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

  tddm_tbt_cordic_f04a48283a: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x11,
      ce_70 => ce_70_sg_x15,
      ch_in => p_ch_out_x2,
      clk_35 => clk_35_sg_x11,
      clk_70 => clk_70_sg_x15,
      din => p_amp_out_x1,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp1/TBT_CORDIC"

entity tbt_cordic_entity_9dc3371de2 is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(24 downto 0);
    q_in: in std_logic_vector(24 downto 0);
    valid_in: in std_logic;
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tddm_tbt_cordic: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x0: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x1: out std_logic_vector(23 downto 0);
    tddm_tbt_cordic_x2: out std_logic_vector(23 downto 0)
  );
end tbt_cordic_entity_9dc3371de2;

architecture structural of tbt_cordic_entity_9dc3371de2 is
  signal ce_35_sg_x12: std_logic;
  signal ce_70_sg_x16: std_logic;
  signal clk_35_sg_x12: std_logic;
  signal clk_70_sg_x16: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal p_amp_out_x2: std_logic_vector(23 downto 0);
  signal p_ch_out_x3: std_logic;
  signal p_phase_out_x1: std_logic_vector(23 downto 0);
  signal phase: std_logic_vector(23 downto 0);
  signal ready: std_logic;
  signal real_x0: std_logic;
  signal register1_q_net_x0: std_logic_vector(24 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register3_q_net_x0: std_logic_vector(24 downto 0);
  signal register6_q_net_x0: std_logic;
  signal reinterpret2_output_port_net: std_logic_vector(23 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(23 downto 0);
  signal valid_out: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x12 <= ce_35;
  ce_70_sg_x16 <= ce_70;
  register2_q_net_x0 <= ch_in;
  clk_35_sg_x12 <= clk_35;
  clk_70_sg_x16 <= clk_70;
  register3_q_net_x0 <= i_in;
  register1_q_net_x0 <= q_in;
  register6_q_net_x0 <= valid_in;
  amp_out <= p_amp_out_x2;
  ch_out <= p_ch_out_x3;
  tddm_tbt_cordic <= down_sample1_q_net_x4;
  tddm_tbt_cordic_x0 <= down_sample2_q_net_x4;
  tddm_tbt_cordic_x1 <= down_sample1_q_net_x5;
  tddm_tbt_cordic_x2 <= down_sample2_q_net_x5;

  rect2pol: entity work.xlcordic_3fb964e2f71602f328fdd11ab57d7304
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      s_axis_cartesian_tdata_imag => register1_q_net_x0,
      s_axis_cartesian_tdata_real => register3_q_net_x0,
      s_axis_cartesian_tuser_user(0) => register2_q_net_x0,
      s_axis_cartesian_tvalid => register6_q_net_x0,
      m_axis_dout_tdata_phase => valid_out,
      m_axis_dout_tdata_real => phase,
      m_axis_dout_tuser_cartesian_tuser(0) => real_x0,
      m_axis_dout_tvalid => ready
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d(0) => real_x0,
      en(0) => ready,
      rst => "0",
      q(0) => p_ch_out_x3
    );

  register4: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => reinterpret2_output_port_net,
      en(0) => ready,
      rst => "0",
      q => p_phase_out_x1
    );

  register5: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x12,
      clk => clk_35_sg_x12,
      d => reinterpret3_output_port_net,
      en(0) => ready,
      rst => "0",
      q => p_amp_out_x2
    );

  reinterpret2: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => valid_out,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_b62f4240f0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => phase,
      output_port => reinterpret3_output_port_net
    );

  tddm_tbt_cordic_9e99bd206d: entity work.tddm_tbt_cordic_entity_9e99bd206d
    port map (
      ce_35 => ce_35_sg_x12,
      ce_70 => ce_70_sg_x16,
      clk_35 => clk_35_sg_x12,
      clk_70 => clk_70_sg_x16,
      tbt_cordic_ch_in => p_ch_out_x3,
      tbt_cordic_din => p_amp_out_x2,
      tbt_cordic_pin => p_phase_out_x1,
      tbt_cordic_ch2_out => down_sample2_q_net_x4,
      tbt_cordic_ch3_out => down_sample1_q_net_x4,
      tbt_cordic_phase0_out => down_sample2_q_net_x5,
      tbt_cordic_phase1_out => down_sample1_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp1/TBT_poly_decim/TDDM_TBT"

entity tddm_tbt_entity_1f4b61e651 is
  port (
    ce_35: in std_logic;
    ce_70: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    tbt_ch_in: in std_logic;
    tbt_i_in: in std_logic_vector(23 downto 0);
    tbt_q_in: in std_logic_vector(23 downto 0);
    poly35_ch2_i_out: out std_logic_vector(23 downto 0);
    poly35_ch2_q_out: out std_logic_vector(23 downto 0);
    poly35_ch3_i_out: out std_logic_vector(23 downto 0);
    poly35_ch3_q_out: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_entity_1f4b61e651;

architecture structural of tddm_tbt_entity_1f4b61e651 is
  signal ce_35_sg_x15: std_logic;
  signal ce_70_sg_x19: std_logic;
  signal clk_35_sg_x15: std_logic;
  signal clk_70_sg_x19: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal register2_q_net_x3: std_logic;
  signal reinterpret_output_port_net_x2: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net_x3: std_logic_vector(23 downto 0);

begin
  ce_35_sg_x15 <= ce_35;
  ce_70_sg_x19 <= ce_70;
  clk_35_sg_x15 <= clk_35;
  clk_70_sg_x19 <= clk_70;
  register2_q_net_x3 <= tbt_ch_in;
  reinterpret_output_port_net_x3 <= tbt_i_in;
  reinterpret_output_port_net_x2 <= tbt_q_in;
  poly35_ch2_i_out <= down_sample2_q_net_x2;
  poly35_ch2_q_out <= down_sample2_q_net_x3;
  poly35_ch3_i_out <= down_sample1_q_net_x2;
  poly35_ch3_q_out <= down_sample1_q_net_x3;

  tddm_tbt_poly_i_b74b709553: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x15,
      ce_70 => ce_70_sg_x19,
      ch_in => register2_q_net_x3,
      clk_35 => clk_35_sg_x15,
      clk_70 => clk_70_sg_x19,
      din => reinterpret_output_port_net_x3,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_tbt_poly_q_4f85d7362a: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x15,
      ce_70 => ce_70_sg_x19,
      ch_in => register2_q_net_x3,
      clk_35 => clk_35_sg_x15,
      clk_70 => clk_70_sg_x19,
      din => reinterpret_output_port_net_x2,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp1/TBT_poly_decim"

entity tbt_poly_decim_entity_bb6f6b5b6a is
  port (
    ce_1: in std_logic;
    ce_35: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    i_out: out std_logic_vector(24 downto 0);
    q_out: out std_logic_vector(24 downto 0);
    tbt_poly_x0: out std_logic;
    tddm_tbt: out std_logic_vector(23 downto 0);
    tddm_tbt_x0: out std_logic_vector(23 downto 0);
    tddm_tbt_x1: out std_logic_vector(23 downto 0);
    tddm_tbt_x2: out std_logic_vector(23 downto 0);
    valid_out: out std_logic
  );
end tbt_poly_decim_entity_bb6f6b5b6a;

architecture structural of tbt_poly_decim_entity_bb6f6b5b6a is
  signal ce_1_sg_x26: std_logic;
  signal ce_35_sg_x16: std_logic;
  signal ce_70_sg_x20: std_logic;
  signal ce_logic_1_sg_x14: std_logic;
  signal clk_1_sg_x26: std_logic;
  signal clk_35_sg_x16: std_logic;
  signal clk_70_sg_x20: std_logic;
  signal down_sample1_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x4: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal register1_q_net_x2: std_logic_vector(24 downto 0);
  signal register2_q_net_x4: std_logic;
  signal register3_q_net_x13: std_logic;
  signal register3_q_net_x2: std_logic_vector(24 downto 0);
  signal register4_q_net_x12: std_logic_vector(23 downto 0);
  signal register5_q_net_x13: std_logic_vector(23 downto 0);
  signal register6_q_net_x1: std_logic;
  signal reinterpret1_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret_output_port_net_x3: std_logic_vector(23 downto 0);
  signal reinterpret_output_port_net_x4: std_logic_vector(23 downto 0);
  signal tbt_poly_event_s_data_chanid_incorrect_net_x0: std_logic;
  signal tbt_poly_m_axis_data_tdata_path0_net: std_logic_vector(24 downto 0);
  signal tbt_poly_m_axis_data_tdata_path1_net: std_logic_vector(24 downto 0);
  signal tbt_poly_m_axis_data_tuser_chanid_net: std_logic;
  signal tbt_poly_m_axis_data_tvalid_net: std_logic;

begin
  ce_1_sg_x26 <= ce_1;
  ce_35_sg_x16 <= ce_35;
  ce_70_sg_x20 <= ce_70;
  ce_logic_1_sg_x14 <= ce_logic_1;
  register3_q_net_x13 <= ch_in;
  clk_1_sg_x26 <= clk_1;
  clk_35_sg_x16 <= clk_35;
  clk_70_sg_x20 <= clk_70;
  register4_q_net_x12 <= i_in;
  register5_q_net_x13 <= q_in;
  ch_out <= register2_q_net_x4;
  i_out <= register3_q_net_x2;
  q_out <= register1_q_net_x2;
  tbt_poly_x0 <= tbt_poly_event_s_data_chanid_incorrect_net_x0;
  tddm_tbt <= down_sample1_q_net_x4;
  tddm_tbt_x0 <= down_sample2_q_net_x4;
  tddm_tbt_x1 <= down_sample1_q_net_x5;
  tddm_tbt_x2 <= down_sample2_q_net_x5;
  valid_out <= register6_q_net_x1;

  register1: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x16,
      clk => clk_35_sg_x16,
      d => reinterpret_output_port_net,
      en(0) => tbt_poly_m_axis_data_tvalid_net,
      rst => "0",
      q => register1_q_net_x2
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x16,
      clk => clk_35_sg_x16,
      d(0) => tbt_poly_m_axis_data_tuser_chanid_net,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x4
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_35_sg_x16,
      clk => clk_35_sg_x16,
      d => reinterpret1_output_port_net,
      en(0) => tbt_poly_m_axis_data_tvalid_net,
      rst => "0",
      q => register3_q_net_x2
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_35_sg_x16,
      clk => clk_35_sg_x16,
      d(0) => tbt_poly_m_axis_data_tvalid_net,
      en => "1",
      rst => "0",
      q(0) => register6_q_net_x1
    );

  reinterpret: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => tbt_poly_m_axis_data_tdata_path1_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => tbt_poly_m_axis_data_tdata_path0_net,
      output_port => reinterpret1_output_port_net
    );

  tbt_poly: entity work.xlfir_compiler_f7093b59b74f3d511e09195b077ec73c
    port map (
      ce => ce_1_sg_x26,
      ce_35 => ce_35_sg_x16,
      ce_logic_1 => ce_logic_1_sg_x14,
      clk => clk_1_sg_x26,
      clk_35 => clk_35_sg_x16,
      clk_logic_1 => clk_1_sg_x26,
      s_axis_data_tdata_path0 => register4_q_net_x12,
      s_axis_data_tdata_path1 => register5_q_net_x13,
      s_axis_data_tuser_chanid(0) => register3_q_net_x13,
      src_ce => ce_1_sg_x26,
      src_clk => clk_1_sg_x26,
      event_s_data_chanid_incorrect => tbt_poly_event_s_data_chanid_incorrect_net_x0,
      m_axis_data_tdata_path0 => tbt_poly_m_axis_data_tdata_path0_net,
      m_axis_data_tdata_path1 => tbt_poly_m_axis_data_tdata_path1_net,
      m_axis_data_tuser_chanid(0) => tbt_poly_m_axis_data_tuser_chanid_net,
      m_axis_data_tvalid => tbt_poly_m_axis_data_tvalid_net
    );

  tddm_tbt_1f4b61e651: entity work.tddm_tbt_entity_1f4b61e651
    port map (
      ce_35 => ce_35_sg_x16,
      ce_70 => ce_70_sg_x20,
      clk_35 => clk_35_sg_x16,
      clk_70 => clk_70_sg_x20,
      tbt_ch_in => register2_q_net_x4,
      tbt_i_in => reinterpret_output_port_net_x4,
      tbt_q_in => reinterpret_output_port_net_x3,
      poly35_ch2_i_out => down_sample2_q_net_x4,
      poly35_ch2_q_out => down_sample2_q_net_x5,
      poly35_ch3_i_out => down_sample1_q_net_x4,
      poly35_ch3_q_out => down_sample1_q_net_x5
    );

  trunc1_c3e3bdeec5: entity work.trunc_entity_e5eda8a5ac
    port map (
      din => register3_q_net_x2,
      dout => reinterpret_output_port_net_x4
    );

  trunc_6a2a4db298: entity work.trunc_entity_e5eda8a5ac
    port map (
      din => register1_q_net_x2,
      dout => reinterpret_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TBT_amp1"

entity tbt_amp1_entity_6e98f85f9f is
  port (
    ce_1: in std_logic;
    ce_35: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ch_in: in std_logic;
    clk_1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in: in std_logic_vector(23 downto 0);
    q_in: in std_logic_vector(23 downto 0);
    amp_out: out std_logic_vector(23 downto 0);
    ch_out: out std_logic;
    tbt_cordic: out std_logic_vector(23 downto 0);
    tbt_cordic_x0: out std_logic_vector(23 downto 0);
    tbt_cordic_x1: out std_logic_vector(23 downto 0);
    tbt_cordic_x2: out std_logic_vector(23 downto 0);
    tbt_poly_decim: out std_logic;
    tbt_poly_decim_x0: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x1: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x2: out std_logic_vector(23 downto 0);
    tbt_poly_decim_x3: out std_logic_vector(23 downto 0)
  );
end tbt_amp1_entity_6e98f85f9f;

architecture structural of tbt_amp1_entity_6e98f85f9f is
  signal ce_1_sg_x27: std_logic;
  signal ce_35_sg_x17: std_logic;
  signal ce_70_sg_x21: std_logic;
  signal ce_logic_1_sg_x15: std_logic;
  signal clk_1_sg_x27: std_logic;
  signal clk_35_sg_x17: std_logic;
  signal clk_70_sg_x21: std_logic;
  signal down_sample1_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x9: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x10: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x11: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x8: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x9: std_logic_vector(23 downto 0);
  signal p_amp_out_x3: std_logic_vector(23 downto 0);
  signal p_ch_out_x4: std_logic;
  signal register1_q_net_x2: std_logic_vector(24 downto 0);
  signal register2_q_net_x4: std_logic;
  signal register3_q_net_x14: std_logic;
  signal register3_q_net_x2: std_logic_vector(24 downto 0);
  signal register4_q_net_x13: std_logic_vector(23 downto 0);
  signal register5_q_net_x14: std_logic_vector(23 downto 0);
  signal register6_q_net_x1: std_logic;
  signal tbt_poly_event_s_data_chanid_incorrect_net_x1: std_logic;

begin
  ce_1_sg_x27 <= ce_1;
  ce_35_sg_x17 <= ce_35;
  ce_70_sg_x21 <= ce_70;
  ce_logic_1_sg_x15 <= ce_logic_1;
  register3_q_net_x14 <= ch_in;
  clk_1_sg_x27 <= clk_1;
  clk_35_sg_x17 <= clk_35;
  clk_70_sg_x21 <= clk_70;
  register4_q_net_x13 <= i_in;
  register5_q_net_x14 <= q_in;
  amp_out <= p_amp_out_x3;
  ch_out <= p_ch_out_x4;
  tbt_cordic <= down_sample1_q_net_x8;
  tbt_cordic_x0 <= down_sample2_q_net_x8;
  tbt_cordic_x1 <= down_sample1_q_net_x9;
  tbt_cordic_x2 <= down_sample2_q_net_x9;
  tbt_poly_decim <= tbt_poly_event_s_data_chanid_incorrect_net_x1;
  tbt_poly_decim_x0 <= down_sample1_q_net_x10;
  tbt_poly_decim_x1 <= down_sample2_q_net_x10;
  tbt_poly_decim_x2 <= down_sample1_q_net_x11;
  tbt_poly_decim_x3 <= down_sample2_q_net_x11;

  tbt_cordic_9dc3371de2: entity work.tbt_cordic_entity_9dc3371de2
    port map (
      ce_35 => ce_35_sg_x17,
      ce_70 => ce_70_sg_x21,
      ch_in => register2_q_net_x4,
      clk_35 => clk_35_sg_x17,
      clk_70 => clk_70_sg_x21,
      i_in => register3_q_net_x2,
      q_in => register1_q_net_x2,
      valid_in => register6_q_net_x1,
      amp_out => p_amp_out_x3,
      ch_out => p_ch_out_x4,
      tddm_tbt_cordic => down_sample1_q_net_x8,
      tddm_tbt_cordic_x0 => down_sample2_q_net_x8,
      tddm_tbt_cordic_x1 => down_sample1_q_net_x9,
      tddm_tbt_cordic_x2 => down_sample2_q_net_x9
    );

  tbt_poly_decim_bb6f6b5b6a: entity work.tbt_poly_decim_entity_bb6f6b5b6a
    port map (
      ce_1 => ce_1_sg_x27,
      ce_35 => ce_35_sg_x17,
      ce_70 => ce_70_sg_x21,
      ce_logic_1 => ce_logic_1_sg_x15,
      ch_in => register3_q_net_x14,
      clk_1 => clk_1_sg_x27,
      clk_35 => clk_35_sg_x17,
      clk_70 => clk_70_sg_x21,
      i_in => register4_q_net_x13,
      q_in => register5_q_net_x14,
      ch_out => register2_q_net_x4,
      i_out => register3_q_net_x2,
      q_out => register1_q_net_x2,
      tbt_poly_x0 => tbt_poly_event_s_data_chanid_incorrect_net_x1,
      tddm_tbt => down_sample1_q_net_x10,
      tddm_tbt_x0 => down_sample2_q_net_x10,
      tddm_tbt_x1 => down_sample1_q_net_x11,
      tddm_tbt_x2 => down_sample2_q_net_x11,
      valid_out => register6_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp/TDDM_tbt_amp_4ch"

entity tddm_tbt_amp_4ch_entity_9f3ac0073e is
  port (
    amp_in0: in std_logic_vector(23 downto 0);
    amp_in1: in std_logic_vector(23 downto 0);
    ce_35: in std_logic;
    ce_70: in std_logic;
    ch_in0: in std_logic;
    ch_in1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    amp_out0: out std_logic_vector(23 downto 0);
    amp_out1: out std_logic_vector(23 downto 0);
    amp_out2: out std_logic_vector(23 downto 0);
    amp_out3: out std_logic_vector(23 downto 0)
  );
end tddm_tbt_amp_4ch_entity_9f3ac0073e;

architecture structural of tddm_tbt_amp_4ch_entity_9f3ac0073e is
  signal ce_35_sg_x20: std_logic;
  signal ce_70_sg_x24: std_logic;
  signal clk_35_sg_x20: std_logic;
  signal clk_70_sg_x24: std_logic;
  signal down_sample1_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x3: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x2: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x3: std_logic_vector(23 downto 0);
  signal p_amp_out_x6: std_logic_vector(23 downto 0);
  signal p_amp_out_x7: std_logic_vector(23 downto 0);
  signal p_ch_out_x7: std_logic;
  signal p_ch_out_x8: std_logic;

begin
  p_amp_out_x6 <= amp_in0;
  p_amp_out_x7 <= amp_in1;
  ce_35_sg_x20 <= ce_35;
  ce_70_sg_x24 <= ce_70;
  p_ch_out_x7 <= ch_in0;
  p_ch_out_x8 <= ch_in1;
  clk_35_sg_x20 <= clk_35;
  clk_70_sg_x24 <= clk_70;
  amp_out0 <= down_sample2_q_net_x2;
  amp_out1 <= down_sample1_q_net_x2;
  amp_out2 <= down_sample2_q_net_x3;
  amp_out3 <= down_sample1_q_net_x3;

  tddm_tbt_amp0_8f2b25894a: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x20,
      ce_70 => ce_70_sg_x24,
      ch_in => p_ch_out_x7,
      clk_35 => clk_35_sg_x20,
      clk_70 => clk_70_sg_x24,
      din => p_amp_out_x6,
      dout_ch0 => down_sample2_q_net_x2,
      dout_ch1 => down_sample1_q_net_x2
    );

  tddm_tbt_amp1_0c4a2e4770: entity work.tddm_tbt_cordic_entity_5b94be40c5
    port map (
      ce_35 => ce_35_sg_x20,
      ce_70 => ce_70_sg_x24,
      ch_in => p_ch_out_x8,
      clk_35 => clk_35_sg_x20,
      clk_70 => clk_70_sg_x24,
      din => p_amp_out_x7,
      dout_ch0 => down_sample2_q_net_x3,
      dout_ch1 => down_sample1_q_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TBT_amp"

entity tbt_amp_entity_cbd277bb0c is
  port (
    ce_1: in std_logic;
    ce_35: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ch_in0: in std_logic;
    ch_in1: in std_logic;
    clk_1: in std_logic;
    clk_35: in std_logic;
    clk_70: in std_logic;
    i_in0: in std_logic_vector(23 downto 0);
    i_in1: in std_logic_vector(23 downto 0);
    q_in0: in std_logic_vector(23 downto 0);
    q_in1: in std_logic_vector(23 downto 0);
    amp_out0: out std_logic_vector(23 downto 0);
    amp_out1: out std_logic_vector(23 downto 0);
    amp_out2: out std_logic_vector(23 downto 0);
    amp_out3: out std_logic_vector(23 downto 0);
    tbt_amp0: out std_logic_vector(23 downto 0);
    tbt_amp0_x0: out std_logic_vector(23 downto 0);
    tbt_amp0_x1: out std_logic_vector(23 downto 0);
    tbt_amp0_x2: out std_logic_vector(23 downto 0);
    tbt_amp0_x3: out std_logic;
    tbt_amp0_x4: out std_logic_vector(23 downto 0);
    tbt_amp0_x5: out std_logic_vector(23 downto 0);
    tbt_amp0_x6: out std_logic_vector(23 downto 0);
    tbt_amp0_x7: out std_logic_vector(23 downto 0);
    tbt_amp1: out std_logic_vector(23 downto 0);
    tbt_amp1_x0: out std_logic_vector(23 downto 0);
    tbt_amp1_x1: out std_logic_vector(23 downto 0);
    tbt_amp1_x2: out std_logic_vector(23 downto 0);
    tbt_amp1_x3: out std_logic;
    tbt_amp1_x4: out std_logic_vector(23 downto 0);
    tbt_amp1_x5: out std_logic_vector(23 downto 0);
    tbt_amp1_x6: out std_logic_vector(23 downto 0);
    tbt_amp1_x7: out std_logic_vector(23 downto 0)
  );
end tbt_amp_entity_cbd277bb0c;

architecture structural of tbt_amp_entity_cbd277bb0c is
  signal ce_1_sg_x28: std_logic;
  signal ce_35_sg_x21: std_logic;
  signal ce_70_sg_x25: std_logic;
  signal ce_logic_1_sg_x16: std_logic;
  signal clk_1_sg_x28: std_logic;
  signal clk_35_sg_x21: std_logic;
  signal clk_70_sg_x25: std_logic;
  signal down_sample1_q_net_x16: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x17: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x19: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x22: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x23: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x24: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x25: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x16: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x17: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x19: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x22: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x23: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x24: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x25: std_logic_vector(23 downto 0);
  signal p_amp_out_x6: std_logic_vector(23 downto 0);
  signal p_amp_out_x7: std_logic_vector(23 downto 0);
  signal p_ch_out_x7: std_logic;
  signal p_ch_out_x8: std_logic;
  signal register3_q_net_x15: std_logic;
  signal register3_q_net_x16: std_logic;
  signal register4_q_net_x14: std_logic_vector(23 downto 0);
  signal register4_q_net_x15: std_logic_vector(23 downto 0);
  signal register5_q_net_x11: std_logic_vector(23 downto 0);
  signal register5_q_net_x15: std_logic_vector(23 downto 0);
  signal tbt_poly_event_s_data_chanid_incorrect_net_x3: std_logic;
  signal tbt_poly_event_s_data_chanid_incorrect_net_x4: std_logic;

begin
  ce_1_sg_x28 <= ce_1;
  ce_35_sg_x21 <= ce_35;
  ce_70_sg_x25 <= ce_70;
  ce_logic_1_sg_x16 <= ce_logic_1;
  register3_q_net_x15 <= ch_in0;
  register3_q_net_x16 <= ch_in1;
  clk_1_sg_x28 <= clk_1;
  clk_35_sg_x21 <= clk_35;
  clk_70_sg_x25 <= clk_70;
  register4_q_net_x14 <= i_in0;
  register4_q_net_x15 <= i_in1;
  register5_q_net_x11 <= q_in0;
  register5_q_net_x15 <= q_in1;
  amp_out0 <= down_sample2_q_net_x24;
  amp_out1 <= down_sample1_q_net_x24;
  amp_out2 <= down_sample2_q_net_x25;
  amp_out3 <= down_sample1_q_net_x25;
  tbt_amp0 <= down_sample1_q_net_x16;
  tbt_amp0_x0 <= down_sample2_q_net_x16;
  tbt_amp0_x1 <= down_sample1_q_net_x17;
  tbt_amp0_x2 <= down_sample2_q_net_x17;
  tbt_amp0_x3 <= tbt_poly_event_s_data_chanid_incorrect_net_x3;
  tbt_amp0_x4 <= down_sample1_q_net_x18;
  tbt_amp0_x5 <= down_sample2_q_net_x18;
  tbt_amp0_x6 <= down_sample1_q_net_x19;
  tbt_amp0_x7 <= down_sample2_q_net_x19;
  tbt_amp1 <= down_sample1_q_net_x20;
  tbt_amp1_x0 <= down_sample2_q_net_x20;
  tbt_amp1_x1 <= down_sample1_q_net_x21;
  tbt_amp1_x2 <= down_sample2_q_net_x21;
  tbt_amp1_x3 <= tbt_poly_event_s_data_chanid_incorrect_net_x4;
  tbt_amp1_x4 <= down_sample1_q_net_x22;
  tbt_amp1_x5 <= down_sample2_q_net_x22;
  tbt_amp1_x6 <= down_sample1_q_net_x23;
  tbt_amp1_x7 <= down_sample2_q_net_x23;

  tbt_amp0_88b1c45f0e: entity work.tbt_amp0_entity_88b1c45f0e
    port map (
      ce_1 => ce_1_sg_x28,
      ce_35 => ce_35_sg_x21,
      ce_70 => ce_70_sg_x25,
      ce_logic_1 => ce_logic_1_sg_x16,
      ch_in => register3_q_net_x15,
      clk_1 => clk_1_sg_x28,
      clk_35 => clk_35_sg_x21,
      clk_70 => clk_70_sg_x25,
      i_in => register4_q_net_x14,
      q_in => register5_q_net_x11,
      amp_out => p_amp_out_x6,
      ch_out => p_ch_out_x7,
      tbt_cordic => down_sample1_q_net_x16,
      tbt_cordic_x0 => down_sample2_q_net_x16,
      tbt_cordic_x1 => down_sample1_q_net_x17,
      tbt_cordic_x2 => down_sample2_q_net_x17,
      tbt_poly_decim => tbt_poly_event_s_data_chanid_incorrect_net_x3,
      tbt_poly_decim_x0 => down_sample1_q_net_x18,
      tbt_poly_decim_x1 => down_sample2_q_net_x18,
      tbt_poly_decim_x2 => down_sample1_q_net_x19,
      tbt_poly_decim_x3 => down_sample2_q_net_x19
    );

  tbt_amp1_6e98f85f9f: entity work.tbt_amp1_entity_6e98f85f9f
    port map (
      ce_1 => ce_1_sg_x28,
      ce_35 => ce_35_sg_x21,
      ce_70 => ce_70_sg_x25,
      ce_logic_1 => ce_logic_1_sg_x16,
      ch_in => register3_q_net_x16,
      clk_1 => clk_1_sg_x28,
      clk_35 => clk_35_sg_x21,
      clk_70 => clk_70_sg_x25,
      i_in => register4_q_net_x15,
      q_in => register5_q_net_x15,
      amp_out => p_amp_out_x7,
      ch_out => p_ch_out_x8,
      tbt_cordic => down_sample1_q_net_x20,
      tbt_cordic_x0 => down_sample2_q_net_x20,
      tbt_cordic_x1 => down_sample1_q_net_x21,
      tbt_cordic_x2 => down_sample2_q_net_x21,
      tbt_poly_decim => tbt_poly_event_s_data_chanid_incorrect_net_x4,
      tbt_poly_decim_x0 => down_sample1_q_net_x22,
      tbt_poly_decim_x1 => down_sample2_q_net_x22,
      tbt_poly_decim_x2 => down_sample1_q_net_x23,
      tbt_poly_decim_x3 => down_sample2_q_net_x23
    );

  tddm_tbt_amp_4ch_9f3ac0073e: entity work.tddm_tbt_amp_4ch_entity_9f3ac0073e
    port map (
      amp_in0 => p_amp_out_x6,
      amp_in1 => p_amp_out_x7,
      ce_35 => ce_35_sg_x21,
      ce_70 => ce_70_sg_x25,
      ch_in0 => p_ch_out_x7,
      ch_in1 => p_ch_out_x8,
      clk_35 => clk_35_sg_x21,
      clk_70 => clk_70_sg_x25,
      amp_out0 => down_sample2_q_net_x24,
      amp_out1 => down_sample1_q_net_x24,
      amp_out2 => down_sample2_q_net_x25,
      amp_out3 => down_sample1_q_net_x25
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_mix/TDM_mix_ch0_1"

entity tdm_mix_ch0_1_entity_b9bb73dd5f is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_logic_1: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    din_ch0: in std_logic_vector(23 downto 0);
    din_ch1: in std_logic_vector(23 downto 0);
    rst: in std_logic;
    ch_out: out std_logic;
    dout: out std_logic_vector(23 downto 0)
  );
end tdm_mix_ch0_1_entity_b9bb73dd5f;

architecture structural of tdm_mix_ch0_1_entity_b9bb73dd5f is
  signal ce_1_sg_x29: std_logic;
  signal ce_2_sg_x31: std_logic;
  signal ce_logic_1_sg_x17: std_logic;
  signal clk_1_sg_x29: std_logic;
  signal clk_2_sg_x31: std_logic;
  signal clock_enable_probe_q_net: std_logic;
  signal constant10_op_net_x0: std_logic;
  signal mux_sel1_op_net: std_logic;
  signal mux_y_net: std_logic_vector(23 downto 0);
  signal register1_q_net_x4: std_logic;
  signal register_q_net_x17: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x8: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x9: std_logic_vector(23 downto 0);
  signal up_sample_ch0_q_net: std_logic_vector(23 downto 0);
  signal up_sample_ch1_q_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x29 <= ce_1;
  ce_2_sg_x31 <= ce_2;
  ce_logic_1_sg_x17 <= ce_logic_1;
  clk_1_sg_x29 <= clk_1;
  clk_2_sg_x31 <= clk_2;
  reinterpret2_output_port_net_x9 <= din_ch0;
  reinterpret2_output_port_net_x8 <= din_ch1;
  constant10_op_net_x0 <= rst;
  ch_out <= register1_q_net_x4;
  dout <= register_q_net_x17;

  clock_enable_probe: entity work.xlceprobe
    generic map (
      d_width => 24,
      q_width => 1
    )
    port map (
      ce => ce_logic_1_sg_x17,
      clk => clk_1_sg_x29,
      d => up_sample_ch0_q_net,
      q(0) => clock_enable_probe_q_net
    );

  mux: entity work.mux_a2121d82da
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => up_sample_ch0_q_net,
      d1 => up_sample_ch1_q_net,
      sel(0) => mux_sel1_op_net,
      y => mux_y_net
    );

  mux_sel1: entity work.counter_41314d726b
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      en(0) => clock_enable_probe_q_net,
      rst(0) => constant10_op_net_x0,
      op(0) => mux_sel1_op_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d(0) => mux_sel1_op_net,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x4
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      d => mux_y_net,
      en => "1",
      rst => "0",
      q => register_q_net_x17
    );

  up_sample_ch0: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => reinterpret2_output_port_net_x9,
      dest_ce => ce_1_sg_x29,
      dest_clk => clk_1_sg_x29,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x31,
      src_clk => clk_2_sg_x31,
      src_clr => '0',
      q => up_sample_ch0_q_net
    );

  up_sample_ch1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => reinterpret2_output_port_net_x8,
      dest_ce => ce_1_sg_x29,
      dest_clk => clk_1_sg_x29,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x31,
      src_clk => clk_2_sg_x31,
      src_clr => '0',
      q => up_sample_ch1_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_mix"

entity tdm_mix_entity_54ce67e6e8 is
  port (
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_logic_1: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    din_ch0: in std_logic_vector(23 downto 0);
    din_ch1: in std_logic_vector(23 downto 0);
    din_ch2: in std_logic_vector(23 downto 0);
    din_ch3: in std_logic_vector(23 downto 0);
    ch_out0: out std_logic;
    ch_out1: out std_logic;
    dout0: out std_logic_vector(23 downto 0);
    dout1: out std_logic_vector(23 downto 0)
  );
end tdm_mix_entity_54ce67e6e8;

architecture structural of tdm_mix_entity_54ce67e6e8 is
  signal ce_1_sg_x31: std_logic;
  signal ce_2_sg_x33: std_logic;
  signal ce_logic_1_sg_x19: std_logic;
  signal clk_1_sg_x31: std_logic;
  signal clk_2_sg_x33: std_logic;
  signal constant10_op_net_x0: std_logic;
  signal constant11_op_net_x0: std_logic;
  signal register1_q_net_x6: std_logic;
  signal register1_q_net_x7: std_logic;
  signal register_q_net_x19: std_logic_vector(23 downto 0);
  signal register_q_net_x20: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x11: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x12: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x13: std_logic_vector(23 downto 0);
  signal reinterpret2_output_port_net_x14: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x31 <= ce_1;
  ce_2_sg_x33 <= ce_2;
  ce_logic_1_sg_x19 <= ce_logic_1;
  clk_1_sg_x31 <= clk_1;
  clk_2_sg_x33 <= clk_2;
  reinterpret2_output_port_net_x14 <= din_ch0;
  reinterpret2_output_port_net_x11 <= din_ch1;
  reinterpret2_output_port_net_x12 <= din_ch2;
  reinterpret2_output_port_net_x13 <= din_ch3;
  ch_out0 <= register1_q_net_x6;
  ch_out1 <= register1_q_net_x7;
  dout0 <= register_q_net_x19;
  dout1 <= register_q_net_x20;

  constant10: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant10_op_net_x0
    );

  constant11: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant11_op_net_x0
    );

  tdm_mix_ch0_1_b9bb73dd5f: entity work.tdm_mix_ch0_1_entity_b9bb73dd5f
    port map (
      ce_1 => ce_1_sg_x31,
      ce_2 => ce_2_sg_x33,
      ce_logic_1 => ce_logic_1_sg_x19,
      clk_1 => clk_1_sg_x31,
      clk_2 => clk_2_sg_x33,
      din_ch0 => reinterpret2_output_port_net_x14,
      din_ch1 => reinterpret2_output_port_net_x11,
      rst => constant10_op_net_x0,
      ch_out => register1_q_net_x6,
      dout => register_q_net_x19
    );

  tdm_mix_ch0_2_e9327141fc: entity work.tdm_mix_ch0_1_entity_b9bb73dd5f
    port map (
      ce_1 => ce_1_sg_x31,
      ce_2 => ce_2_sg_x33,
      ce_logic_1 => ce_logic_1_sg_x19,
      clk_1 => clk_1_sg_x31,
      clk_2 => clk_2_sg_x33,
      din_ch0 => reinterpret2_output_port_net_x12,
      din_ch1 => reinterpret2_output_port_net_x13,
      rst => constant11_op_net_x0,
      ch_out => register1_q_net_x7,
      dout => register_q_net_x20
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_monit"

entity tdm_monit_entity_6e38292ecb is
  port (
    ce_1: in std_logic;
    ce_2240: in std_logic;
    ce_560: in std_logic;
    ce_logic_560: in std_logic;
    clk_1: in std_logic;
    clk_2240: in std_logic;
    clk_560: in std_logic;
    din_ch0: in std_logic_vector(23 downto 0);
    din_ch1: in std_logic_vector(23 downto 0);
    din_ch2: in std_logic_vector(23 downto 0);
    din_ch3: in std_logic_vector(23 downto 0);
    rst: in std_logic;
    ch_out: out std_logic_vector(1 downto 0);
    dout: out std_logic_vector(23 downto 0)
  );
end tdm_monit_entity_6e38292ecb;

architecture structural of tdm_monit_entity_6e38292ecb is
  signal ce_1_sg_x32: std_logic;
  signal ce_2240_sg_x26: std_logic;
  signal ce_560_sg_x2: std_logic;
  signal ce_logic_560_sg_x2: std_logic;
  signal ch_out_x2: std_logic_vector(1 downto 0);
  signal clk_1_sg_x32: std_logic;
  signal clk_2240_sg_x26: std_logic;
  signal clk_560_sg_x2: std_logic;
  signal clock_enable_probe_q_net: std_logic;
  signal constant10_op_net_x0: std_logic;
  signal dout_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x19: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x18: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x19: std_logic_vector(23 downto 0);
  signal mux_sel_op_net: std_logic_vector(1 downto 0);
  signal mux_y_net: std_logic_vector(23 downto 0);
  signal up_sample_ch0_q_net: std_logic_vector(23 downto 0);
  signal up_sample_ch1_q_net: std_logic_vector(23 downto 0);
  signal up_sample_ch2_q_net: std_logic_vector(23 downto 0);
  signal up_sample_ch3_q_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x32 <= ce_1;
  ce_2240_sg_x26 <= ce_2240;
  ce_560_sg_x2 <= ce_560;
  ce_logic_560_sg_x2 <= ce_logic_560;
  clk_1_sg_x32 <= clk_1;
  clk_2240_sg_x26 <= clk_2240;
  clk_560_sg_x2 <= clk_560;
  down_sample2_q_net_x18 <= din_ch0;
  down_sample1_q_net_x18 <= din_ch1;
  down_sample2_q_net_x19 <= din_ch2;
  down_sample1_q_net_x19 <= din_ch3;
  constant10_op_net_x0 <= rst;
  ch_out <= ch_out_x2;
  dout <= dout_x2;

  clock_enable_probe: entity work.xlceprobe
    generic map (
      d_width => 24,
      q_width => 1
    )
    port map (
      ce => ce_logic_560_sg_x2,
      clk => clk_560_sg_x2,
      d => up_sample_ch0_q_net,
      q(0) => clock_enable_probe_q_net
    );

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 2,
      ds_ratio => 560,
      latency => 1,
      phase => 559,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 2
    )
    port map (
      d => mux_sel_op_net,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x32,
      src_clk => clk_1_sg_x32,
      src_clr => '0',
      q => ch_out_x2
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      ds_ratio => 560,
      latency => 1,
      phase => 559,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => mux_y_net,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x32,
      src_clk => clk_1_sg_x32,
      src_clr => '0',
      q => dout_x2
    );

  mux: entity work.mux_f062741975
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => up_sample_ch0_q_net,
      d1 => up_sample_ch1_q_net,
      d2 => up_sample_ch2_q_net,
      d3 => up_sample_ch3_q_net,
      sel => mux_sel_op_net,
      y => mux_y_net
    );

  mux_sel: entity work.xlcounter_free
    generic map (
      core_name0 => "cntr_11_0_eb46eda57512a5a4",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      en(0) => clock_enable_probe_q_net,
      rst(0) => constant10_op_net_x0,
      op => mux_sel_op_net
    );

  up_sample_ch0: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => down_sample2_q_net_x18,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x26,
      src_clk => clk_2240_sg_x26,
      src_clr => '0',
      q => up_sample_ch0_q_net
    );

  up_sample_ch1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => down_sample1_q_net_x18,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x26,
      src_clk => clk_2240_sg_x26,
      src_clr => '0',
      q => up_sample_ch1_q_net
    );

  up_sample_ch2: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => down_sample2_q_net_x19,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x26,
      src_clk => clk_2240_sg_x26,
      src_clr => '0',
      q => up_sample_ch2_q_net
    );

  up_sample_ch3: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 24,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 24
    )
    port map (
      d => down_sample1_q_net_x19,
      dest_ce => ce_560_sg_x2,
      dest_clk => clk_560_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x26,
      src_clk => clk_2240_sg_x26,
      src_clr => '0',
      q => up_sample_ch3_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_monit_1/downsample"

entity downsample_entity_f33f90217c is
  port (
    ce_1: in std_logic;
    ce_2500: in std_logic;
    ce_5600000: in std_logic;
    clk_1: in std_logic;
    clk_2500: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(1 downto 0);
    dout: out std_logic_vector(1 downto 0)
  );
end downsample_entity_f33f90217c;

architecture structural of downsample_entity_f33f90217c is
  signal ce_1_sg_x33: std_logic;
  signal ce_2500_sg_x0: std_logic;
  signal ce_5600000_sg_x8: std_logic;
  signal clk_1_sg_x33: std_logic;
  signal clk_2500_sg_x0: std_logic;
  signal clk_5600000_sg_x8: std_logic;
  signal down_sample5_q_net: std_logic_vector(1 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(1 downto 0);
  signal mux_sel_op_net_x0: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x33 <= ce_1;
  ce_2500_sg_x0 <= ce_2500;
  ce_5600000_sg_x8 <= ce_5600000;
  clk_1_sg_x33 <= clk_1;
  clk_2500_sg_x0 <= clk_2500;
  clk_5600000_sg_x8 <= clk_5600000;
  mux_sel_op_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 2,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 2
    )
    port map (
      d => down_sample5_q_net,
      dest_ce => ce_5600000_sg_x8,
      dest_clk => clk_5600000_sg_x8,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2500_sg_x0,
      src_clk => clk_2500_sg_x0,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 2,
      ds_ratio => 2500,
      latency => 1,
      phase => 2499,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 2
    )
    port map (
      d => mux_sel_op_net_x0,
      dest_ce => ce_2500_sg_x0,
      dest_clk => clk_2500_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x33,
      src_clk => clk_1_sg_x33,
      src_clr => '0',
      q => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_monit_1/downsample1"

entity downsample1_entity_312d531c6b is
  port (
    ce_1: in std_logic;
    ce_2500: in std_logic;
    ce_5600000: in std_logic;
    clk_1: in std_logic;
    clk_2500: in std_logic;
    clk_5600000: in std_logic;
    din: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(25 downto 0)
  );
end downsample1_entity_312d531c6b;

architecture structural of downsample1_entity_312d531c6b is
  signal ce_1_sg_x34: std_logic;
  signal ce_2500_sg_x1: std_logic;
  signal ce_5600000_sg_x9: std_logic;
  signal clk_1_sg_x34: std_logic;
  signal clk_2500_sg_x1: std_logic;
  signal clk_5600000_sg_x9: std_logic;
  signal down_sample5_q_net: std_logic_vector(25 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(25 downto 0);
  signal mux_y_net_x0: std_logic_vector(25 downto 0);

begin
  ce_1_sg_x34 <= ce_1;
  ce_2500_sg_x1 <= ce_2500;
  ce_5600000_sg_x9 <= ce_5600000;
  clk_1_sg_x34 <= clk_1;
  clk_2500_sg_x1 <= clk_2500;
  clk_5600000_sg_x9 <= clk_5600000;
  mux_y_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => down_sample5_q_net,
      dest_ce => ce_5600000_sg_x9,
      dest_clk => clk_5600000_sg_x9,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2500_sg_x1,
      src_clk => clk_2500_sg_x1,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 2500,
      latency => 1,
      phase => 2499,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => mux_y_net_x0,
      dest_ce => ce_2500_sg_x1,
      dest_clk => clk_2500_sg_x1,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x34,
      src_clk => clk_1_sg_x34,
      src_clr => '0',
      q => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/TDM_monit_1"

entity tdm_monit_1_entity_746ecf54b0 is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_2500: in std_logic;
    ce_5600000: in std_logic;
    ce_logic_5600000: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_2500: in std_logic;
    clk_5600000: in std_logic;
    din_ch0: in std_logic_vector(25 downto 0);
    din_ch1: in std_logic_vector(25 downto 0);
    din_ch2: in std_logic_vector(25 downto 0);
    din_ch3: in std_logic_vector(25 downto 0);
    rst: in std_logic;
    ch_out: out std_logic_vector(1 downto 0);
    dout: out std_logic_vector(25 downto 0)
  );
end tdm_monit_1_entity_746ecf54b0;

architecture structural of tdm_monit_1_entity_746ecf54b0 is
  signal ce_1_sg_x35: std_logic;
  signal ce_22400000_sg_x10: std_logic;
  signal ce_2500_sg_x2: std_logic;
  signal ce_5600000_sg_x10: std_logic;
  signal ce_logic_5600000_sg_x0: std_logic;
  signal clk_1_sg_x35: std_logic;
  signal clk_22400000_sg_x10: std_logic;
  signal clk_2500_sg_x2: std_logic;
  signal clk_5600000_sg_x10: std_logic;
  signal clock_enable_probe_q_net: std_logic;
  signal concat1_y_net_x0: std_logic_vector(25 downto 0);
  signal concat2_y_net_x0: std_logic_vector(25 downto 0);
  signal concat3_y_net_x0: std_logic_vector(25 downto 0);
  signal concat_y_net_x0: std_logic_vector(25 downto 0);
  signal constant11_op_net_x0: std_logic;
  signal down_sample_q_net_x2: std_logic_vector(1 downto 0);
  signal down_sample_q_net_x3: std_logic_vector(25 downto 0);
  signal mux_sel_op_net_x0: std_logic_vector(1 downto 0);
  signal mux_y_net_x0: std_logic_vector(25 downto 0);
  signal up_sample_ch0_q_net: std_logic_vector(25 downto 0);
  signal up_sample_ch1_q_net: std_logic_vector(25 downto 0);
  signal up_sample_ch2_q_net: std_logic_vector(25 downto 0);
  signal up_sample_ch3_q_net: std_logic_vector(25 downto 0);

begin
  ce_1_sg_x35 <= ce_1;
  ce_22400000_sg_x10 <= ce_22400000;
  ce_2500_sg_x2 <= ce_2500;
  ce_5600000_sg_x10 <= ce_5600000;
  ce_logic_5600000_sg_x0 <= ce_logic_5600000;
  clk_1_sg_x35 <= clk_1;
  clk_22400000_sg_x10 <= clk_22400000;
  clk_2500_sg_x2 <= clk_2500;
  clk_5600000_sg_x10 <= clk_5600000;
  concat_y_net_x0 <= din_ch0;
  concat1_y_net_x0 <= din_ch1;
  concat2_y_net_x0 <= din_ch2;
  concat3_y_net_x0 <= din_ch3;
  constant11_op_net_x0 <= rst;
  ch_out <= down_sample_q_net_x2;
  dout <= down_sample_q_net_x3;

  clock_enable_probe: entity work.xlceprobe
    generic map (
      d_width => 26,
      q_width => 1
    )
    port map (
      ce => ce_logic_5600000_sg_x0,
      clk => clk_5600000_sg_x10,
      d => up_sample_ch0_q_net,
      q(0) => clock_enable_probe_q_net
    );

  downsample1_312d531c6b: entity work.downsample1_entity_312d531c6b
    port map (
      ce_1 => ce_1_sg_x35,
      ce_2500 => ce_2500_sg_x2,
      ce_5600000 => ce_5600000_sg_x10,
      clk_1 => clk_1_sg_x35,
      clk_2500 => clk_2500_sg_x2,
      clk_5600000 => clk_5600000_sg_x10,
      din => mux_y_net_x0,
      dout => down_sample_q_net_x3
    );

  downsample_f33f90217c: entity work.downsample_entity_f33f90217c
    port map (
      ce_1 => ce_1_sg_x35,
      ce_2500 => ce_2500_sg_x2,
      ce_5600000 => ce_5600000_sg_x10,
      clk_1 => clk_1_sg_x35,
      clk_2500 => clk_2500_sg_x2,
      clk_5600000 => clk_5600000_sg_x10,
      din => mux_sel_op_net_x0,
      dout => down_sample_q_net_x2
    );

  mux: entity work.mux_187c900130
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => up_sample_ch0_q_net,
      d1 => up_sample_ch1_q_net,
      d2 => up_sample_ch2_q_net,
      d3 => up_sample_ch3_q_net,
      sel => mux_sel_op_net_x0,
      y => mux_y_net_x0
    );

  mux_sel: entity work.xlcounter_free
    generic map (
      core_name0 => "cntr_11_0_eb46eda57512a5a4",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x35,
      clk => clk_1_sg_x35,
      clr => '0',
      en(0) => clock_enable_probe_q_net,
      rst(0) => constant11_op_net_x0,
      op => mux_sel_op_net_x0
    );

  up_sample_ch0: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => concat_y_net_x0,
      dest_ce => ce_5600000_sg_x10,
      dest_clk => clk_5600000_sg_x10,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x10,
      src_clk => clk_22400000_sg_x10,
      src_clr => '0',
      q => up_sample_ch0_q_net
    );

  up_sample_ch1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => concat1_y_net_x0,
      dest_ce => ce_5600000_sg_x10,
      dest_clk => clk_5600000_sg_x10,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x10,
      src_clk => clk_22400000_sg_x10,
      src_clr => '0',
      q => up_sample_ch1_q_net
    );

  up_sample_ch2: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => concat2_y_net_x0,
      dest_ce => ce_5600000_sg_x10,
      dest_clk => clk_5600000_sg_x10,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x10,
      src_clk => clk_22400000_sg_x10,
      src_clr => '0',
      q => up_sample_ch2_q_net
    );

  up_sample_ch3: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => concat3_y_net_x0,
      dest_ce => ce_5600000_sg_x10,
      dest_clk => clk_5600000_sg_x10,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x10,
      src_clk => clk_22400000_sg_x10,
      src_clr => '0',
      q => up_sample_ch3_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/convert_filt"

entity convert_filt_entity_fda412c1bf is
  port (
    din: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(24 downto 0)
  );
end convert_filt_entity_fda412c1bf;

architecture structural of convert_filt_entity_fda412c1bf is
  signal down_sample_q_net_x4: std_logic_vector(25 downto 0);
  signal extractor1_dout_net: std_logic_vector(24 downto 0);
  signal reinterpret5_output_port_net_x0: std_logic_vector(24 downto 0);

begin
  down_sample_q_net_x4 <= din;
  dout <= reinterpret5_output_port_net_x0;

  extractor1: entity work.bitbasher_a756ba0096
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      din => down_sample_q_net_x4,
      dout => extractor1_dout_net
    );

  reinterpret5: entity work.reinterpret_60ea556961
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => extractor1_dout_net,
      output_port => reinterpret5_output_port_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb/DataReg_En"

entity datareg_en_entity_79473f9ed1 is
  port (
    ce_1: in std_logic;
    clk_1: in std_logic;
    din: in std_logic_vector(24 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(24 downto 0);
    valid: out std_logic
  );
end datareg_en_entity_79473f9ed1;

architecture structural of datareg_en_entity_79473f9ed1 is
  signal ce_1_sg_x36: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal divider_dout_valid_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x36 <= ce_1;
  clk_1_sg_x36 <= clk_1;
  reinterpret1_output_port_net_x0 <= din;
  divider_dout_valid_x0 <= en;
  dout <= register_q_net_x0;
  valid <= register1_q_net_x0;

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => divider_dout_valid_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d => reinterpret1_output_port_net_x0,
      en(0) => divider_dout_valid_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb/DataReg_En3"

entity datareg_en3_entity_6643090018 is
  port (
    ce_1: in std_logic;
    clk_1: in std_logic;
    din: in std_logic_vector(24 downto 0);
    en: in std_logic;
    dout: out std_logic_vector(24 downto 0);
    valid: out std_logic
  );
end datareg_en3_entity_6643090018;

architecture structural of datareg_en3_entity_6643090018 is
  signal ce_1_sg_x39: std_logic;
  signal clk_1_sg_x39: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal delay1_q_net_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x39 <= ce_1;
  clk_1_sg_x39 <= clk_1;
  convert_dout_net_x0 <= din;
  delay1_q_net_x0 <= en;
  dout <= register_q_net_x0;
  valid <= register1_q_net_x0;

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      d(0) => delay1_q_net_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x39,
      clk => clk_1_sg_x39,
      d => convert_dout_net_x0,
      en(0) => delay1_q_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb/pulse_stretcher"

entity pulse_stretcher_entity_9893378b63 is
  port (
    ce_1: in std_logic;
    clk_1: in std_logic;
    clr: in std_logic;
    pulse_in: in std_logic;
    extd_out: out std_logic
  );
end pulse_stretcher_entity_9893378b63;

architecture structural of pulse_stretcher_entity_9893378b63 is
  signal ce_1_sg_x40: std_logic;
  signal ce_70_x0: std_logic;
  signal clk_1_sg_x40: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal register1_q_net_x1: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x40 <= ce_1;
  clk_1_sg_x40 <= clk_1;
  ce_70_x0 <= clr;
  register1_q_net_x1 <= pulse_in;
  extd_out <= logical3_y_net_x0;

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      clr => '0',
      ip(0) => ce_70_x0,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register_q_net,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register1_q_net_x1,
      d1(0) => logical1_y_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register1_q_net_x1,
      d1(0) => register_q_net,
      y(0) => logical3_y_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      d(0) => logical2_y_net,
      en => "1",
      rst => "0",
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_fofb"

entity delta_sigma_fofb_entity_ee61e649ea is
  port (
    a: in std_logic_vector(23 downto 0);
    b: in std_logic_vector(23 downto 0);
    c: in std_logic_vector(23 downto 0);
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_2240: in std_logic;
    ce_logic_2240: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    clk_2240: in std_logic;
    d: in std_logic_vector(23 downto 0);
    ds_thres: in std_logic_vector(25 downto 0);
    q: out std_logic_vector(24 downto 0);
    q_valid: out std_logic;
    sum_valid: out std_logic;
    sum_x0: out std_logic_vector(24 downto 0);
    x: out std_logic_vector(24 downto 0);
    x_valid: out std_logic;
    y: out std_logic_vector(24 downto 0);
    y_valid: out std_logic
  );
end delta_sigma_fofb_entity_ee61e649ea;

architecture structural of delta_sigma_fofb_entity_ee61e649ea is
  signal a_plus_b_s_net: std_logic_vector(24 downto 0);
  signal a_plus_c_s_net: std_logic_vector(24 downto 0);
  signal a_plus_d_s_net: std_logic_vector(24 downto 0);
  signal assert10_dout_net_x1: std_logic;
  signal assert11_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x1: std_logic;
  signal assert1_dout_net_x0: std_logic;
  signal assert5_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert6_dout_net_x0: std_logic;
  signal assert8_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert9_dout_net_x1: std_logic;
  signal assert_dout_net: std_logic;
  signal b_plus_c_s_net: std_logic_vector(24 downto 0);
  signal b_plus_d_s_net: std_logic_vector(24 downto 0);
  signal c_plus_d_s_net: std_logic_vector(24 downto 0);
  signal ce_1_sg_x48: std_logic;
  signal ce_2240_sg_x27: std_logic;
  signal ce_2_sg_x34: std_logic;
  signal ce_70_x3: std_logic;
  signal ce_logic_2240_sg_x0: std_logic;
  signal clk_1_sg_x48: std_logic;
  signal clk_2240_sg_x27: std_logic;
  signal clk_2_sg_x34: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal del_sig_div_fofb_thres_i_net_x0: std_logic_vector(25 downto 0);
  signal delay1_q_net_x0: std_logic;
  signal delay_q_net: std_logic_vector(25 downto 0);
  signal delta_q_s_net: std_logic_vector(25 downto 0);
  signal delta_x_s_net: std_logic_vector(25 downto 0);
  signal delta_y_s_net: std_logic_vector(25 downto 0);
  signal din: std_logic_vector(25 downto 0);
  signal dividend_data: std_logic_vector(25 downto 0);
  signal dividend_ready: std_logic;
  signal dividend_ready_x0: std_logic;
  signal dividend_valid_x0: std_logic;
  signal dividend_valid_x1: std_logic;
  signal dividend_valid_x2: std_logic;
  signal divider_dout_fracc: std_logic_vector(24 downto 0);
  signal divider_dout_valid_x0: std_logic;
  signal divisor_data: std_logic_vector(25 downto 0);
  signal divisor_data_x0: std_logic_vector(25 downto 0);
  signal divisor_ready: std_logic;
  signal divisor_valid_x0: std_logic;
  signal dout_down_x1: std_logic_vector(24 downto 0);
  signal dout_stretch: std_logic_vector(24 downto 0);
  signal down_sample1_q_net: std_logic_vector(24 downto 0);
  signal down_sample1_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample2_q_net: std_logic;
  signal down_sample2_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample3_q_net: std_logic_vector(24 downto 0);
  signal down_sample4_q_net: std_logic;
  signal down_sample5_q_net: std_logic_vector(24 downto 0);
  signal down_sample6_q_net: std_logic;
  signal down_sample7_q_net: std_logic_vector(24 downto 0);
  signal down_sample8_q_net: std_logic;
  signal down_sample_q_net: std_logic_vector(25 downto 0);
  signal expression1_dout_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical3_y_net_x2: std_logic;
  signal logical3_y_net_x3: std_logic;
  signal logical3_y_net_x4: std_logic;
  signal logical3_y_net_x5: std_logic;
  signal logical3_y_net_x6: std_logic;
  signal logical3_y_net_x7: std_logic;
  signal q_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal q_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal q_divider_s_axis_dividend_tready_net: std_logic;
  signal q_divider_s_axis_divisor_tready_net: std_logic;
  signal re_x0: std_logic;
  signal re_x1: std_logic;
  signal register10_q_net: std_logic_vector(25 downto 0);
  signal register11_q_net: std_logic_vector(24 downto 0);
  signal register12_q_net: std_logic_vector(24 downto 0);
  signal register13_q_net: std_logic_vector(24 downto 0);
  signal register14_q_net: std_logic_vector(25 downto 0);
  signal register1_q_net: std_logic_vector(24 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register1_q_net_x2: std_logic;
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x4: std_logic;
  signal register2_q_net: std_logic_vector(24 downto 0);
  signal register3_q_net: std_logic_vector(24 downto 0);
  signal register4_q_net: std_logic_vector(24 downto 0);
  signal register5_q_net: std_logic_vector(24 downto 0);
  signal register6_q_net: std_logic_vector(24 downto 0);
  signal register7_q_net: std_logic_vector(25 downto 0);
  signal register_q_net_x0: std_logic_vector(24 downto 0);
  signal register_q_net_x1: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal register_q_net_x3: std_logic_vector(24 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret7_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret8_output_port_net: std_logic_vector(25 downto 0);
  signal relational_op_net: std_logic;
  signal sum_s_net: std_logic_vector(25 downto 0);
  signal up_sample2_q_net: std_logic_vector(25 downto 0);
  signal up_sample4_q_net: std_logic_vector(25 downto 0);
  signal up_sample6_q_net: std_logic_vector(25 downto 0);
  signal up_sample_q_net: std_logic_vector(25 downto 0);
  signal valid_ds_down_x1: std_logic;
  signal x_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal x_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal x_divider_s_axis_divisor_tready_net: std_logic;

begin
  down_sample2_q_net_x20 <= a;
  down_sample1_q_net_x20 <= b;
  down_sample2_q_net_x21 <= c;
  ce_1_sg_x48 <= ce_1;
  ce_2_sg_x34 <= ce_2;
  ce_2240_sg_x27 <= ce_2240;
  ce_logic_2240_sg_x0 <= ce_logic_2240;
  clk_1_sg_x48 <= clk_1;
  clk_2_sg_x34 <= clk_2;
  clk_2240_sg_x27 <= clk_2240;
  down_sample1_q_net_x21 <= d;
  del_sig_div_fofb_thres_i_net_x0 <= ds_thres;
  q <= assert8_dout_net_x1;
  q_valid <= assert9_dout_net_x1;
  sum_valid <= assert12_dout_net_x1;
  sum_x0 <= assert11_dout_net_x1;
  x <= assert5_dout_net_x1;
  x_valid <= assert10_dout_net_x1;
  y <= dout_down_x1;
  y_valid <= valid_ds_down_x1;

  a_plus_b: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x20,
      b => down_sample1_q_net_x20,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_b_s_net
    );

  a_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x20,
      b => down_sample2_q_net_x21,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_c_s_net
    );

  a_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x20,
      b => down_sample1_q_net_x21,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_d_s_net
    );

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => q_divider_s_axis_dividend_tready_net,
      dout(0) => assert1_dout_net_x0
    );

  assert10: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample6_q_net,
      dout(0) => assert10_dout_net_x1
    );

  assert11: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample7_q_net,
      dout => assert11_dout_net_x1
    );

  assert12: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample8_q_net,
      dout(0) => assert12_dout_net_x1
    );

  assert2: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready_x0,
      dout(0) => re_x0
    );

  assert3: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready,
      dout(0) => re_x1
    );

  assert4: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample1_q_net,
      dout => dout_down_x1
    );

  assert5: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample5_q_net,
      dout => assert5_dout_net_x1
    );

  assert6: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => expression1_dout_net,
      dout(0) => assert6_dout_net_x0
    );

  assert7: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample2_q_net,
      dout(0) => valid_ds_down_x1
    );

  assert8: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample3_q_net,
      dout => assert8_dout_net_x1
    );

  assert9: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample4_q_net,
      dout(0) => assert9_dout_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => relational_op_net,
      dout(0) => assert_dout_net
    );

  b_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x20,
      b => down_sample2_q_net_x21,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => b_plus_c_s_net
    );

  b_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x20,
      b => down_sample1_q_net_x21,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => b_plus_d_s_net
    );

  c_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x21,
      b => down_sample1_q_net_x21,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => c_plus_d_s_net
    );

  ce1: entity work.xlceprobe
    generic map (
      d_width => 1,
      q_width => 1
    )
    port map (
      ce => ce_logic_2240_sg_x0,
      clk => clk_2240_sg_x27,
      d(0) => assert_dout_net,
      q(0) => ce_70_x3
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 22,
      din_width => 26,
      dout_arith => 2,
      dout_bin_pt => 21,
      dout_width => 25,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlRound
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      clr => '0',
      din => delay_q_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  datareg_en1_3225c09afc: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      din => reinterpret2_output_port_net_x0,
      en => q_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x1,
      valid => register1_q_net_x2
    );

  datareg_en2_5b5f4b61b7: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      din => reinterpret3_output_port_net_x0,
      en => x_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x2,
      valid => register1_q_net_x3
    );

  datareg_en3_6643090018: entity work.datareg_en3_entity_6643090018
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      din => convert_dout_net_x0,
      en => delay1_q_net_x0,
      dout => register_q_net_x3,
      valid => register1_q_net_x4
    );

  datareg_en_79473f9ed1: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      din => reinterpret1_output_port_net_x0,
      en => divider_dout_valid_x0,
      dout => register_q_net_x0,
      valid => register1_q_net_x1
    );

  delay: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 26
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d => reinterpret8_output_port_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d(0) => logical3_y_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  delta_q: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register5_q_net,
      b => register6_q_net,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => delta_q_s_net
    );

  delta_x: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register1_q_net,
      b => register3_q_net,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => delta_x_s_net
    );

  delta_y: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register2_q_net,
      b => register4_q_net,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => delta_y_s_net
    );

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      ds_ratio => 1120,
      latency => 1,
      phase => 1119,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register14_q_net,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x34,
      src_clk => clk_2_sg_x34,
      src_clr => '0',
      q => down_sample_q_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => dout_stretch,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample1_q_net
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x0,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q(0) => down_sample2_q_net
    );

  down_sample3: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => register11_q_net,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample3_q_net
    );

  down_sample4: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x1,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q(0) => down_sample4_q_net
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => register12_q_net,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample5_q_net
    );

  down_sample6: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x2,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q(0) => down_sample6_q_net
    );

  down_sample7: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 25,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 25
    )
    port map (
      d => register13_q_net,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q => down_sample7_q_net
    );

  down_sample8: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 2240,
      latency => 1,
      phase => 2239,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x3,
      dest_ce => ce_2240_sg_x27,
      dest_clk => clk_2240_sg_x27,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x48,
      src_clk => clk_1_sg_x48,
      src_clr => '0',
      q(0) => down_sample8_q_net
    );

  expression1: entity work.expr_375d7bbece
    port map (
      a(0) => x_divider_s_axis_divisor_tready_net,
      b(0) => divisor_ready,
      c(0) => q_divider_s_axis_divisor_tready_net,
      ce => '0',
      clk => '0',
      clr => '0',
      dout(0) => expression1_dout_net
    );

  pulse_stretcher1_f6401a1a3d: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x2,
      extd_out => logical3_y_net_x1
    );

  pulse_stretcher2_38948aaba0: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x3,
      extd_out => logical3_y_net_x2
    );

  pulse_stretcher3_816d954034: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x4,
      extd_out => logical3_y_net_x3
    );

  pulse_stretcher4_5d505b900f: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => assert6_dout_net_x0,
      pulse_in => divisor_valid_x0,
      extd_out => logical3_y_net_x4
    );

  pulse_stretcher5_bee4540339: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => re_x0,
      pulse_in => dividend_valid_x0,
      extd_out => logical3_y_net_x5
    );

  pulse_stretcher6_f82d879b1c: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => assert1_dout_net_x0,
      pulse_in => dividend_valid_x1,
      extd_out => logical3_y_net_x6
    );

  pulse_stretcher7_2406c4a105: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => re_x1,
      pulse_in => dividend_valid_x2,
      extd_out => logical3_y_net_x7
    );

  pulse_stretcher_9893378b63: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x48,
      clk_1 => clk_1_sg_x48,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x1,
      extd_out => logical3_y_net_x0
    );

  q_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      s_axis_dividend_tdata_dividend => reinterpret7_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x6,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => q_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => q_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => q_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => q_divider_s_axis_divisor_tready_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => b_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register10: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => delta_q_s_net,
      en => "1",
      rst => "0",
      q => register10_q_net
    );

  register11: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d => register_q_net_x1,
      en => "1",
      rst => "0",
      q => register11_q_net
    );

  register12: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d => register_q_net_x2,
      en => "1",
      rst => "0",
      q => register12_q_net
    );

  register13: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d => register_q_net_x3,
      en => "1",
      rst => "0",
      q => register13_q_net
    );

  register14: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x34,
      clk => clk_2_sg_x34,
      d => del_sig_div_fofb_thres_i_net_x0,
      en => "1",
      rst => "0",
      q => register14_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => a_plus_b_s_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => a_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => c_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => a_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => b_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register6_q_net
    );

  register7: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => delta_x_s_net,
      en => "1",
      rst => "0",
      q => register7_q_net
    );

  register8: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => sum_s_net,
      en => "1",
      rst => "0",
      q => divisor_data
    );

  register9: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      d => delta_y_s_net,
      en => "1",
      rst => "0",
      q => din
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      d => register_q_net_x0,
      en => "1",
      rst => "0",
      q => dout_stretch
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divider_dout_fracc,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => q_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => x_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample6_q_net,
      output_port => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample2_q_net,
      output_port => divisor_data_x0
    );

  reinterpret6: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample_q_net,
      output_port => dividend_data
    );

  reinterpret7: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample4_q_net,
      output_port => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divisor_data_x0,
      output_port => reinterpret8_output_port_net
    );

  relational: entity work.relational_416cfcae1e
    port map (
      a => divisor_data,
      b => down_sample_q_net,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      op(0) => relational_op_net
    );

  sum: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_3537d66a2361cd1e",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register3_q_net,
      b => register1_q_net,
      ce => ce_2240_sg_x27,
      clk => clk_2240_sg_x27,
      clr => '0',
      en => "1",
      s => sum_s_net
    );

  up_sample: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => din,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q => up_sample_q_net
    );

  up_sample1: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q(0) => dividend_valid_x0
    );

  up_sample2: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => divisor_data,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q => up_sample2_q_net
    );

  up_sample3: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q(0) => divisor_valid_x0
    );

  up_sample4: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register10_q_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q => up_sample4_q_net
    );

  up_sample5: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q(0) => dividend_valid_x1
    );

  up_sample6: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register7_q_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q => up_sample6_q_net
    );

  up_sample7: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x48,
      dest_clk => clk_1_sg_x48,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2240_sg_x27,
      src_clk => clk_2240_sg_x27,
      src_clr => '0',
      q(0) => dividend_valid_x2
    );

  x_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      s_axis_dividend_tdata_dividend => reinterpret4_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x7,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => x_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => x_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => dividend_ready,
      s_axis_divisor_tready => x_divider_s_axis_divisor_tready_net
    );

  y_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x48,
      clk => clk_1_sg_x48,
      s_axis_dividend_tdata_dividend => dividend_data,
      s_axis_dividend_tvalid => logical3_y_net_x5,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => divider_dout_fracc,
      m_axis_dout_tvalid => divider_dout_valid_x0,
      s_axis_dividend_tready => dividend_ready_x0,
      s_axis_divisor_tready => divisor_ready
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/downsample1"

entity downsample1_entity_4c88924603 is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_5000: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_5000: in std_logic;
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(24 downto 0)
  );
end downsample1_entity_4c88924603;

architecture structural of downsample1_entity_4c88924603 is
  signal ce_1_sg_x53: std_logic;
  signal ce_22400000_sg_x11: std_logic;
  signal ce_5000_sg_x0: std_logic;
  signal clk_1_sg_x53: std_logic;
  signal clk_22400000_sg_x11: std_logic;
  signal clk_5000_sg_x0: std_logic;
  signal down_sample5_q_net: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(24 downto 0);
  signal register13_q_net_x0: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x53 <= ce_1;
  ce_22400000_sg_x11 <= ce_22400000;
  ce_5000_sg_x0 <= ce_5000;
  clk_1_sg_x53 <= clk_1;
  clk_22400000_sg_x11 <= clk_22400000;
  clk_5000_sg_x0 <= clk_5000;
  register13_q_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 25,
      ds_ratio => 4480,
      latency => 1,
      phase => 4479,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 25
    )
    port map (
      d => down_sample5_q_net,
      dest_ce => ce_22400000_sg_x11,
      dest_clk => clk_22400000_sg_x11,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5000_sg_x0,
      src_clk => clk_5000_sg_x0,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 25,
      ds_ratio => 5000,
      latency => 1,
      phase => 4999,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 25
    )
    port map (
      d => register13_q_net_x0,
      dest_ce => ce_5000_sg_x0,
      dest_clk => clk_5000_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x53,
      src_clk => clk_1_sg_x53,
      src_clr => '0',
      q => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/downsample2"

entity downsample2_entity_891f07b1a7 is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_5000: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_5000: in std_logic;
    din: in std_logic;
    dout: out std_logic
  );
end downsample2_entity_891f07b1a7;

architecture structural of downsample2_entity_891f07b1a7 is
  signal ce_1_sg_x54: std_logic;
  signal ce_22400000_sg_x12: std_logic;
  signal ce_5000_sg_x1: std_logic;
  signal clk_1_sg_x54: std_logic;
  signal clk_22400000_sg_x12: std_logic;
  signal clk_5000_sg_x1: std_logic;
  signal down_sample5_q_net: std_logic;
  signal down_sample_q_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;

begin
  ce_1_sg_x54 <= ce_1;
  ce_22400000_sg_x12 <= ce_22400000;
  ce_5000_sg_x1 <= ce_5000;
  clk_1_sg_x54 <= clk_1;
  clk_22400000_sg_x12 <= clk_22400000;
  clk_5000_sg_x1 <= clk_5000;
  logical3_y_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 4480,
      latency => 1,
      phase => 4479,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => down_sample5_q_net,
      dest_ce => ce_22400000_sg_x12,
      dest_clk => clk_22400000_sg_x12,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5000_sg_x1,
      src_clk => clk_5000_sg_x1,
      src_clr => '0',
      q(0) => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 5000,
      latency => 1,
      phase => 4999,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x0,
      dest_ce => ce_5000_sg_x1,
      dest_clk => clk_5000_sg_x1,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x54,
      src_clk => clk_1_sg_x54,
      src_clr => '0',
      q(0) => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/downsample3"

entity downsample3_entity_dba589aaee is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_5000: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_5000: in std_logic;
    din: in std_logic_vector(24 downto 0);
    dout: out std_logic_vector(24 downto 0)
  );
end downsample3_entity_dba589aaee;

architecture structural of downsample3_entity_dba589aaee is
  signal ce_1_sg_x55: std_logic;
  signal ce_22400000_sg_x13: std_logic;
  signal ce_5000_sg_x2: std_logic;
  signal clk_1_sg_x55: std_logic;
  signal clk_22400000_sg_x13: std_logic;
  signal clk_5000_sg_x2: std_logic;
  signal down_sample5_q_net: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(24 downto 0);
  signal register12_q_net_x0: std_logic_vector(24 downto 0);

begin
  ce_1_sg_x55 <= ce_1;
  ce_22400000_sg_x13 <= ce_22400000;
  ce_5000_sg_x2 <= ce_5000;
  clk_1_sg_x55 <= clk_1;
  clk_22400000_sg_x13 <= clk_22400000;
  clk_5000_sg_x2 <= clk_5000;
  register12_q_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 4480,
      latency => 1,
      phase => 4479,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => down_sample5_q_net,
      dest_ce => ce_22400000_sg_x13,
      dest_clk => clk_22400000_sg_x13,
      dest_clr => '0',
      en => "1",
      src_ce => ce_5000_sg_x2,
      src_clk => clk_5000_sg_x2,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 5000,
      latency => 1,
      phase => 4999,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => register12_q_net_x0,
      dest_ce => ce_5000_sg_x2,
      dest_clk => clk_5000_sg_x2,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x55,
      src_clk => clk_1_sg_x55,
      src_clr => '0',
      q => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/downsample7"

entity downsample7_entity_b85055cb62 is
  port (
    ce_10000: in std_logic;
    ce_2: in std_logic;
    ce_44800000: in std_logic;
    clk_10000: in std_logic;
    clk_2: in std_logic;
    clk_44800000: in std_logic;
    din: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(25 downto 0)
  );
end downsample7_entity_b85055cb62;

architecture structural of downsample7_entity_b85055cb62 is
  signal ce_10000_sg_x0: std_logic;
  signal ce_2_sg_x35: std_logic;
  signal ce_44800000_sg_x0: std_logic;
  signal clk_10000_sg_x0: std_logic;
  signal clk_2_sg_x35: std_logic;
  signal clk_44800000_sg_x0: std_logic;
  signal down_sample5_q_net: std_logic_vector(25 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(25 downto 0);
  signal register14_q_net_x0: std_logic_vector(25 downto 0);

begin
  ce_10000_sg_x0 <= ce_10000;
  ce_2_sg_x35 <= ce_2;
  ce_44800000_sg_x0 <= ce_44800000;
  clk_10000_sg_x0 <= clk_10000;
  clk_2_sg_x35 <= clk_2;
  clk_44800000_sg_x0 <= clk_44800000;
  register14_q_net_x0 <= din;
  dout <= down_sample_q_net_x0;

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      ds_ratio => 4480,
      latency => 1,
      phase => 4479,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => down_sample5_q_net,
      dest_ce => ce_44800000_sg_x0,
      dest_clk => clk_44800000_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_10000_sg_x0,
      src_clk => clk_10000_sg_x0,
      src_clr => '0',
      q => down_sample_q_net_x0
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      ds_ratio => 5000,
      latency => 1,
      phase => 4999,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register14_q_net_x0,
      dest_ce => ce_10000_sg_x0,
      dest_clk => clk_10000_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x35,
      src_clk => clk_2_sg_x35,
      src_clr => '0',
      q => down_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/upsample_copy_pad"

entity upsample_copy_pad_entity_86c97eac4f is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_4480: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_4480: in std_logic;
    din: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(25 downto 0)
  );
end upsample_copy_pad_entity_86c97eac4f;

architecture structural of upsample_copy_pad_entity_86c97eac4f is
  signal ce_1_sg_x69: std_logic;
  signal ce_22400000_sg_x19: std_logic;
  signal ce_4480_sg_x0: std_logic;
  signal clk_1_sg_x69: std_logic;
  signal clk_22400000_sg_x19: std_logic;
  signal clk_4480_sg_x0: std_logic;
  signal register10_q_net_x0: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x0: std_logic_vector(25 downto 0);
  signal up_sample5_q_net: std_logic_vector(25 downto 0);

begin
  ce_1_sg_x69 <= ce_1;
  ce_22400000_sg_x19 <= ce_22400000;
  ce_4480_sg_x0 <= ce_4480;
  clk_1_sg_x69 <= clk_1;
  clk_22400000_sg_x19 <= clk_22400000;
  clk_4480_sg_x0 <= clk_4480;
  register10_q_net_x0 <= din;
  dout <= up_sample1_q_net_x0;

  up_sample1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => up_sample5_q_net,
      dest_ce => ce_1_sg_x69,
      dest_clk => clk_1_sg_x69,
      dest_clr => '0',
      en => "1",
      src_ce => ce_4480_sg_x0,
      src_clk => clk_4480_sg_x0,
      src_clr => '0',
      q => up_sample1_q_net_x0
    );

  up_sample5: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register10_q_net_x0,
      dest_ce => ce_4480_sg_x0,
      dest_clk => clk_4480_sg_x0,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x19,
      src_clk => clk_22400000_sg_x19,
      src_clr => '0',
      q => up_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/upsample_copy_pad1"

entity upsample_copy_pad1_entity_edde199d79 is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_4480: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_4480: in std_logic;
    din_x0: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(25 downto 0)
  );
end upsample_copy_pad1_entity_edde199d79;

architecture structural of upsample_copy_pad1_entity_edde199d79 is
  signal ce_1_sg_x70: std_logic;
  signal ce_22400000_sg_x20: std_logic;
  signal ce_4480_sg_x1: std_logic;
  signal clk_1_sg_x70: std_logic;
  signal clk_22400000_sg_x20: std_logic;
  signal clk_4480_sg_x1: std_logic;
  signal din_x1: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x0: std_logic_vector(25 downto 0);
  signal up_sample5_q_net: std_logic_vector(25 downto 0);

begin
  ce_1_sg_x70 <= ce_1;
  ce_22400000_sg_x20 <= ce_22400000;
  ce_4480_sg_x1 <= ce_4480;
  clk_1_sg_x70 <= clk_1;
  clk_22400000_sg_x20 <= clk_22400000;
  clk_4480_sg_x1 <= clk_4480;
  din_x1 <= din_x0;
  dout <= up_sample1_q_net_x0;

  up_sample1: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => up_sample5_q_net,
      dest_ce => ce_1_sg_x70,
      dest_clk => clk_1_sg_x70,
      dest_clr => '0',
      en => "1",
      src_ce => ce_4480_sg_x1,
      src_clk => clk_4480_sg_x1,
      src_clr => '0',
      q => up_sample1_q_net_x0
    );

  up_sample5: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => din_x1,
      dest_ce => ce_4480_sg_x1,
      dest_clk => clk_4480_sg_x1,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x20,
      src_clk => clk_22400000_sg_x20,
      src_clr => '0',
      q => up_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit/upsample_zero_pad"

entity upsample_zero_pad_entity_e334b63be9 is
  port (
    ce_1: in std_logic;
    ce_22400000: in std_logic;
    ce_4480: in std_logic;
    clk_1: in std_logic;
    clk_22400000: in std_logic;
    clk_4480: in std_logic;
    din: in std_logic;
    dout: out std_logic
  );
end upsample_zero_pad_entity_e334b63be9;

architecture structural of upsample_zero_pad_entity_e334b63be9 is
  signal assert13_dout_net_x0: std_logic;
  signal ce_1_sg_x73: std_logic;
  signal ce_22400000_sg_x23: std_logic;
  signal ce_4480_sg_x4: std_logic;
  signal clk_1_sg_x73: std_logic;
  signal clk_22400000_sg_x23: std_logic;
  signal clk_4480_sg_x4: std_logic;
  signal up_sample1_q_net_x1: std_logic;
  signal up_sample5_q_net: std_logic;

begin
  ce_1_sg_x73 <= ce_1;
  ce_22400000_sg_x23 <= ce_22400000;
  ce_4480_sg_x4 <= ce_4480;
  clk_1_sg_x73 <= clk_1;
  clk_22400000_sg_x23 <= clk_22400000;
  clk_4480_sg_x4 <= clk_4480;
  assert13_dout_net_x0 <= din;
  dout <= up_sample1_q_net_x1;

  up_sample1: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => up_sample5_q_net,
      dest_ce => ce_1_sg_x73,
      dest_clk => clk_1_sg_x73,
      dest_clr => '0',
      en => "1",
      src_ce => ce_4480_sg_x4,
      src_clk => clk_4480_sg_x4,
      src_clr => '0',
      q(0) => up_sample1_q_net_x1
    );

  up_sample5: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert13_dout_net_x0,
      dest_ce => ce_4480_sg_x4,
      dest_clk => clk_4480_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_22400000_sg_x23,
      src_clk => clk_22400000_sg_x23,
      src_clr => '0',
      q(0) => up_sample5_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_monit"

entity delta_sigma_monit_entity_a8f8b81626 is
  port (
    a: in std_logic_vector(23 downto 0);
    b: in std_logic_vector(23 downto 0);
    c: in std_logic_vector(23 downto 0);
    ce_1: in std_logic;
    ce_10000: in std_logic;
    ce_2: in std_logic;
    ce_22400000: in std_logic;
    ce_4480: in std_logic;
    ce_44800000: in std_logic;
    ce_5000: in std_logic;
    ce_logic_22400000: in std_logic;
    clk_1: in std_logic;
    clk_10000: in std_logic;
    clk_2: in std_logic;
    clk_22400000: in std_logic;
    clk_4480: in std_logic;
    clk_44800000: in std_logic;
    clk_5000: in std_logic;
    d: in std_logic_vector(23 downto 0);
    ds_thres: in std_logic_vector(25 downto 0);
    q: out std_logic_vector(24 downto 0);
    q_valid: out std_logic;
    sum_valid: out std_logic;
    sum_x0: out std_logic_vector(24 downto 0);
    x: out std_logic_vector(24 downto 0);
    x_valid: out std_logic;
    y: out std_logic_vector(24 downto 0);
    y_valid: out std_logic
  );
end delta_sigma_monit_entity_a8f8b81626;

architecture structural of delta_sigma_monit_entity_a8f8b81626 is
  signal a_plus_b_s_net: std_logic_vector(24 downto 0);
  signal a_plus_c_s_net: std_logic_vector(24 downto 0);
  signal a_plus_d_s_net: std_logic_vector(24 downto 0);
  signal assert10_dout_net_x1: std_logic;
  signal assert11_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x1: std_logic;
  signal assert13_dout_net_x3: std_logic;
  signal assert2_dout_net_x0: std_logic;
  signal assert4_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert5_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert6_dout_net_x0: std_logic;
  signal assert9_dout_net_x1: std_logic;
  signal b_plus_c_s_net: std_logic_vector(24 downto 0);
  signal b_plus_d_s_net: std_logic_vector(24 downto 0);
  signal c_plus_d_s_net: std_logic_vector(24 downto 0);
  signal ce_10000_sg_x1: std_logic;
  signal ce_1_sg_x77: std_logic;
  signal ce_22400000_sg_x27: std_logic;
  signal ce_2_sg_x36: std_logic;
  signal ce_44800000_sg_x1: std_logic;
  signal ce_4480_sg_x8: std_logic;
  signal ce_5000_sg_x8: std_logic;
  signal ce_70_x3: std_logic;
  signal ce_logic_22400000_sg_x0: std_logic;
  signal clk_10000_sg_x1: std_logic;
  signal clk_1_sg_x77: std_logic;
  signal clk_22400000_sg_x27: std_logic;
  signal clk_2_sg_x36: std_logic;
  signal clk_44800000_sg_x1: std_logic;
  signal clk_4480_sg_x8: std_logic;
  signal clk_5000_sg_x8: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal del_sig_div_monit_thres_i_net_x0: std_logic_vector(25 downto 0);
  signal delay1_q_net_x0: std_logic;
  signal delay_q_net: std_logic_vector(25 downto 0);
  signal delta_q_s_net: std_logic_vector(25 downto 0);
  signal delta_x_s_net: std_logic_vector(25 downto 0);
  signal delta_y_s_net: std_logic_vector(25 downto 0);
  signal din_x1: std_logic_vector(25 downto 0);
  signal dividend_data: std_logic_vector(25 downto 0);
  signal dividend_ready: std_logic;
  signal dividend_ready_x0: std_logic;
  signal divider_dout_fracc: std_logic_vector(24 downto 0);
  signal divider_dout_valid_x0: std_logic;
  signal divisor_data: std_logic_vector(25 downto 0);
  signal divisor_data_x0: std_logic_vector(25 downto 0);
  signal divisor_ready: std_logic;
  signal dout_down_x1: std_logic_vector(24 downto 0);
  signal dout_stretch_x0: std_logic_vector(24 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample_q_net_x0: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x1: std_logic;
  signal down_sample_q_net_x2: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x3: std_logic;
  signal down_sample_q_net_x4: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x5: std_logic;
  signal down_sample_q_net_x6: std_logic_vector(25 downto 0);
  signal down_sample_q_net_x7: std_logic_vector(24 downto 0);
  signal down_sample_q_net_x8: std_logic;
  signal expression1_dout_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical3_y_net_x2: std_logic;
  signal logical3_y_net_x3: std_logic;
  signal logical3_y_net_x4: std_logic;
  signal logical3_y_net_x5: std_logic;
  signal logical3_y_net_x6: std_logic;
  signal logical3_y_net_x7: std_logic;
  signal q_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal q_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal q_divider_s_axis_dividend_tready_net: std_logic;
  signal q_divider_s_axis_divisor_tready_net: std_logic;
  signal re_x0: std_logic;
  signal re_x1: std_logic;
  signal register10_q_net_x0: std_logic_vector(25 downto 0);
  signal register11_q_net_x0: std_logic_vector(24 downto 0);
  signal register12_q_net_x0: std_logic_vector(24 downto 0);
  signal register13_q_net_x0: std_logic_vector(24 downto 0);
  signal register14_q_net_x0: std_logic_vector(25 downto 0);
  signal register1_q_net: std_logic_vector(24 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register1_q_net_x2: std_logic;
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x4: std_logic;
  signal register2_q_net: std_logic_vector(24 downto 0);
  signal register3_q_net: std_logic_vector(24 downto 0);
  signal register4_q_net: std_logic_vector(24 downto 0);
  signal register5_q_net: std_logic_vector(24 downto 0);
  signal register6_q_net: std_logic_vector(24 downto 0);
  signal register7_q_net_x0: std_logic_vector(25 downto 0);
  signal register_q_net_x0: std_logic_vector(24 downto 0);
  signal register_q_net_x1: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal register_q_net_x3: std_logic_vector(24 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret7_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret8_output_port_net: std_logic_vector(25 downto 0);
  signal relational_op_net: std_logic;
  signal sum_s_net: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x0: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x1: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x2: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x3: std_logic_vector(25 downto 0);
  signal up_sample1_q_net_x4: std_logic;
  signal up_sample1_q_net_x5: std_logic;
  signal up_sample1_q_net_x6: std_logic;
  signal up_sample1_q_net_x7: std_logic;
  signal valid_ds_down_x1: std_logic;
  signal x_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal x_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal x_divider_s_axis_divisor_tready_net: std_logic;

begin
  down_sample2_q_net_x5 <= a;
  down_sample1_q_net_x5 <= b;
  down_sample3_q_net_x5 <= c;
  ce_1_sg_x77 <= ce_1;
  ce_10000_sg_x1 <= ce_10000;
  ce_2_sg_x36 <= ce_2;
  ce_22400000_sg_x27 <= ce_22400000;
  ce_4480_sg_x8 <= ce_4480;
  ce_44800000_sg_x1 <= ce_44800000;
  ce_5000_sg_x8 <= ce_5000;
  ce_logic_22400000_sg_x0 <= ce_logic_22400000;
  clk_1_sg_x77 <= clk_1;
  clk_10000_sg_x1 <= clk_10000;
  clk_2_sg_x36 <= clk_2;
  clk_22400000_sg_x27 <= clk_22400000;
  clk_4480_sg_x8 <= clk_4480;
  clk_44800000_sg_x1 <= clk_44800000;
  clk_5000_sg_x8 <= clk_5000;
  down_sample4_q_net_x5 <= d;
  del_sig_div_monit_thres_i_net_x0 <= ds_thres;
  q <= assert4_dout_net_x1;
  q_valid <= assert9_dout_net_x1;
  sum_valid <= assert10_dout_net_x1;
  sum_x0 <= assert5_dout_net_x1;
  x <= assert11_dout_net_x1;
  x_valid <= assert12_dout_net_x1;
  y <= dout_down_x1;
  y_valid <= valid_ds_down_x1;

  a_plus_b: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x5,
      b => down_sample1_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_b_s_net
    );

  a_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x5,
      b => down_sample3_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_c_s_net
    );

  a_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x5,
      b => down_sample4_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => a_plus_d_s_net
    );

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready_x0,
      dout(0) => re_x0
    );

  assert10: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample_q_net_x1,
      dout(0) => assert10_dout_net_x1
    );

  assert11: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample_q_net_x2,
      dout => assert11_dout_net_x1
    );

  assert12: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample_q_net_x3,
      dout(0) => assert12_dout_net_x1
    );

  assert13: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => relational_op_net,
      dout(0) => assert13_dout_net_x3
    );

  assert2: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => q_divider_s_axis_dividend_tready_net,
      dout(0) => assert2_dout_net_x0
    );

  assert3: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready,
      dout(0) => re_x1
    );

  assert4: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample_q_net_x7,
      dout => assert4_dout_net_x1
    );

  assert5: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample_q_net_x0,
      dout => assert5_dout_net_x1
    );

  assert6: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => expression1_dout_net,
      dout(0) => assert6_dout_net_x0
    );

  assert7: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample_q_net_x4,
      dout => dout_down_x1
    );

  assert8: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample_q_net_x5,
      dout(0) => valid_ds_down_x1
    );

  assert9: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample_q_net_x8,
      dout(0) => assert9_dout_net_x1
    );

  b_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x5,
      b => down_sample3_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => b_plus_c_s_net
    );

  b_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x5,
      b => down_sample4_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => b_plus_d_s_net
    );

  c_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample3_q_net_x5,
      b => down_sample4_q_net_x5,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => c_plus_d_s_net
    );

  ce1: entity work.xlceprobe
    generic map (
      d_width => 1,
      q_width => 1
    )
    port map (
      ce => ce_logic_22400000_sg_x0,
      clk => clk_22400000_sg_x27,
      d(0) => assert13_dout_net_x3,
      q(0) => ce_70_x3
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 22,
      din_width => 26,
      dout_arith => 2,
      dout_bin_pt => 21,
      dout_width => 25,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlRound
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      din => delay_q_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  datareg_en1_0658df0e73: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      din => reinterpret2_output_port_net_x0,
      en => q_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x1,
      valid => register1_q_net_x2
    );

  datareg_en2_b216d22f41: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      din => reinterpret3_output_port_net_x0,
      en => x_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x2,
      valid => register1_q_net_x3
    );

  datareg_en3_352b935ccb: entity work.datareg_en3_entity_6643090018
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      din => convert_dout_net_x0,
      en => delay1_q_net_x0,
      dout => register_q_net_x3,
      valid => register1_q_net_x4
    );

  datareg_en_8be792d5b9: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      din => reinterpret1_output_port_net_x0,
      en => divider_dout_valid_x0,
      dout => register_q_net_x0,
      valid => register1_q_net_x1
    );

  delay: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 26
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d => reinterpret8_output_port_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => logical3_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  delta_q: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register5_q_net,
      b => register6_q_net,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => delta_q_s_net
    );

  delta_x: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register1_q_net,
      b => register3_q_net,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => delta_x_s_net
    );

  delta_y: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register2_q_net,
      b => register4_q_net,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => delta_y_s_net
    );

  downsample1_4c88924603: entity work.downsample1_entity_4c88924603
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => register13_q_net_x0,
      dout => down_sample_q_net_x0
    );

  downsample2_891f07b1a7: entity work.downsample2_entity_891f07b1a7
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => logical3_y_net_x4,
      dout => down_sample_q_net_x1
    );

  downsample3_dba589aaee: entity work.downsample3_entity_dba589aaee
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => register12_q_net_x0,
      dout => down_sample_q_net_x2
    );

  downsample4_c9912c17cb: entity work.downsample2_entity_891f07b1a7
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => logical3_y_net_x3,
      dout => down_sample_q_net_x3
    );

  downsample5_5d411d5dea: entity work.downsample3_entity_dba589aaee
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => dout_stretch_x0,
      dout => down_sample_q_net_x4
    );

  downsample6_d7e68015e5: entity work.downsample2_entity_891f07b1a7
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => logical3_y_net_x1,
      dout => down_sample_q_net_x5
    );

  downsample7_b85055cb62: entity work.downsample7_entity_b85055cb62
    port map (
      ce_10000 => ce_10000_sg_x1,
      ce_2 => ce_2_sg_x36,
      ce_44800000 => ce_44800000_sg_x1,
      clk_10000 => clk_10000_sg_x1,
      clk_2 => clk_2_sg_x36,
      clk_44800000 => clk_44800000_sg_x1,
      din => register14_q_net_x0,
      dout => down_sample_q_net_x6
    );

  downsample8_69d7284f0d: entity work.downsample3_entity_dba589aaee
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => register11_q_net_x0,
      dout => down_sample_q_net_x7
    );

  downsample9_f5ac9b8db2: entity work.downsample2_entity_891f07b1a7
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_5000 => ce_5000_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_5000 => clk_5000_sg_x8,
      din => logical3_y_net_x2,
      dout => down_sample_q_net_x8
    );

  expression1: entity work.expr_375d7bbece
    port map (
      a(0) => x_divider_s_axis_divisor_tready_net,
      b(0) => divisor_ready,
      c(0) => q_divider_s_axis_divisor_tready_net,
      ce => '0',
      clk => '0',
      clr => '0',
      dout(0) => expression1_dout_net
    );

  pulse_stretcher1_427f70e3c7: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x2,
      extd_out => logical3_y_net_x2
    );

  pulse_stretcher2_9a61283281: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x3,
      extd_out => logical3_y_net_x3
    );

  pulse_stretcher3_864c3e16a6: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x4,
      extd_out => logical3_y_net_x4
    );

  pulse_stretcher4_8dfd1c8928: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => assert6_dout_net_x0,
      pulse_in => up_sample1_q_net_x6,
      extd_out => logical3_y_net_x0
    );

  pulse_stretcher5_ac376595d0: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => re_x0,
      pulse_in => up_sample1_q_net_x5,
      extd_out => logical3_y_net_x5
    );

  pulse_stretcher6_694b81e6b2: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => assert2_dout_net_x0,
      pulse_in => up_sample1_q_net_x4,
      extd_out => logical3_y_net_x6
    );

  pulse_stretcher7_bb8174efbd: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => re_x1,
      pulse_in => up_sample1_q_net_x7,
      extd_out => logical3_y_net_x7
    );

  pulse_stretcher_6bf297451d: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x77,
      clk_1 => clk_1_sg_x77,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x1,
      extd_out => logical3_y_net_x1
    );

  q_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      s_axis_dividend_tdata_dividend => reinterpret7_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x6,
      s_axis_divisor_tdata_divisor => divisor_data,
      s_axis_divisor_tvalid => logical3_y_net_x0,
      m_axis_dout_tdata_fractional => q_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => q_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => q_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => q_divider_s_axis_divisor_tready_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => b_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register10: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => delta_q_s_net,
      en => "1",
      rst => "0",
      q => register10_q_net_x0
    );

  register11: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d => register_q_net_x1,
      en => "1",
      rst => "0",
      q => register11_q_net_x0
    );

  register12: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d => register_q_net_x2,
      en => "1",
      rst => "0",
      q => register12_q_net_x0
    );

  register13: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d => register_q_net_x3,
      en => "1",
      rst => "0",
      q => register13_q_net_x0
    );

  register14: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x36,
      clk => clk_2_sg_x36,
      d => del_sig_div_monit_thres_i_net_x0,
      en => "1",
      rst => "0",
      q => register14_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => a_plus_b_s_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => a_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => c_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => a_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => b_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register6_q_net
    );

  register7: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => delta_x_s_net,
      en => "1",
      rst => "0",
      q => register7_q_net_x0
    );

  register8: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => sum_s_net,
      en => "1",
      rst => "0",
      q => divisor_data_x0
    );

  register9: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      d => delta_y_s_net,
      en => "1",
      rst => "0",
      q => din_x1
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d => register_q_net_x0,
      en => "1",
      rst => "0",
      q => dout_stretch_x0
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divider_dout_fracc,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => q_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => x_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample1_q_net_x3,
      output_port => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample1_q_net_x2,
      output_port => divisor_data
    );

  reinterpret6: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample1_q_net_x1,
      output_port => dividend_data
    );

  reinterpret7: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample1_q_net_x0,
      output_port => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divisor_data,
      output_port => reinterpret8_output_port_net
    );

  relational: entity work.relational_416cfcae1e
    port map (
      a => divisor_data_x0,
      b => down_sample_q_net_x6,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      op(0) => relational_op_net
    );

  sum: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_3537d66a2361cd1e",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register3_q_net,
      b => register1_q_net,
      ce => ce_22400000_sg_x27,
      clk => clk_22400000_sg_x27,
      clr => '0',
      en => "1",
      s => sum_s_net
    );

  upsample_copy_pad1_edde199d79: entity work.upsample_copy_pad1_entity_edde199d79
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din_x0 => din_x1,
      dout => up_sample1_q_net_x1
    );

  upsample_copy_pad2_46599e345b: entity work.upsample_copy_pad_entity_86c97eac4f
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => divisor_data_x0,
      dout => up_sample1_q_net_x2
    );

  upsample_copy_pad3_3571daa38f: entity work.upsample_copy_pad_entity_86c97eac4f
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => register7_q_net_x0,
      dout => up_sample1_q_net_x3
    );

  upsample_copy_pad_86c97eac4f: entity work.upsample_copy_pad_entity_86c97eac4f
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => register10_q_net_x0,
      dout => up_sample1_q_net_x0
    );

  upsample_zero_pad1_2044d1ec3f: entity work.upsample_zero_pad_entity_e334b63be9
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => assert13_dout_net_x3,
      dout => up_sample1_q_net_x5
    );

  upsample_zero_pad2_7f2f8f8620: entity work.upsample_zero_pad_entity_e334b63be9
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => assert13_dout_net_x3,
      dout => up_sample1_q_net_x6
    );

  upsample_zero_pad3_f0b4acbf28: entity work.upsample_zero_pad_entity_e334b63be9
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => assert13_dout_net_x3,
      dout => up_sample1_q_net_x7
    );

  upsample_zero_pad_e334b63be9: entity work.upsample_zero_pad_entity_e334b63be9
    port map (
      ce_1 => ce_1_sg_x77,
      ce_22400000 => ce_22400000_sg_x27,
      ce_4480 => ce_4480_sg_x8,
      clk_1 => clk_1_sg_x77,
      clk_22400000 => clk_22400000_sg_x27,
      clk_4480 => clk_4480_sg_x8,
      din => assert13_dout_net_x3,
      dout => up_sample1_q_net_x4
    );

  x_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      s_axis_dividend_tdata_dividend => reinterpret4_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x7,
      s_axis_divisor_tdata_divisor => divisor_data,
      s_axis_divisor_tvalid => logical3_y_net_x0,
      m_axis_dout_tdata_fractional => x_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => x_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => dividend_ready,
      s_axis_divisor_tready => x_divider_s_axis_divisor_tready_net
    );

  y_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      s_axis_dividend_tdata_dividend => dividend_data,
      s_axis_dividend_tvalid => logical3_y_net_x5,
      s_axis_divisor_tdata_divisor => divisor_data,
      s_axis_divisor_tvalid => logical3_y_net_x0,
      m_axis_dout_tdata_fractional => divider_dout_fracc,
      m_axis_dout_tvalid => divider_dout_valid_x0,
      s_axis_dividend_tready => dividend_ready_x0,
      s_axis_divisor_tready => divisor_ready
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/delta-sigma_tbt"

entity delta_sigma_tbt_entity_bbfa8a8a69 is
  port (
    a: in std_logic_vector(23 downto 0);
    b: in std_logic_vector(23 downto 0);
    c: in std_logic_vector(23 downto 0);
    ce_1: in std_logic;
    ce_2: in std_logic;
    ce_70: in std_logic;
    ce_logic_70: in std_logic;
    clk_1: in std_logic;
    clk_2: in std_logic;
    clk_70: in std_logic;
    d: in std_logic_vector(23 downto 0);
    ds_thres: in std_logic_vector(25 downto 0);
    q: out std_logic_vector(24 downto 0);
    q_valid: out std_logic;
    sum_valid: out std_logic;
    sum_x0: out std_logic_vector(24 downto 0);
    x: out std_logic_vector(24 downto 0);
    x_valid: out std_logic;
    y: out std_logic_vector(24 downto 0);
    y_valid: out std_logic
  );
end delta_sigma_tbt_entity_bbfa8a8a69;

architecture structural of delta_sigma_tbt_entity_bbfa8a8a69 is
  signal a_plus_b_s_net: std_logic_vector(24 downto 0);
  signal a_plus_c_s_net: std_logic_vector(24 downto 0);
  signal a_plus_d_s_net: std_logic_vector(24 downto 0);
  signal assert10_dout_net_x1: std_logic;
  signal assert11_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x1: std_logic;
  signal assert1_dout_net_x0: std_logic;
  signal assert5_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert6_dout_net_x0: std_logic;
  signal assert8_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert9_dout_net_x1: std_logic;
  signal assert_dout_net: std_logic;
  signal b_plus_c_s_net: std_logic_vector(24 downto 0);
  signal b_plus_d_s_net: std_logic_vector(24 downto 0);
  signal c_plus_d_s_net: std_logic_vector(24 downto 0);
  signal ce_1_sg_x90: std_logic;
  signal ce_2_sg_x37: std_logic;
  signal ce_70_sg_x26: std_logic;
  signal ce_70_x3: std_logic;
  signal ce_logic_70_sg_x0: std_logic;
  signal clk_1_sg_x90: std_logic;
  signal clk_2_sg_x37: std_logic;
  signal clk_70_sg_x26: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal del_sig_div_tbt_thres_i_net_x0: std_logic_vector(25 downto 0);
  signal delay1_q_net_x0: std_logic;
  signal delay_q_net: std_logic_vector(25 downto 0);
  signal delta_q_s_net: std_logic_vector(25 downto 0);
  signal delta_x_s_net: std_logic_vector(25 downto 0);
  signal delta_y_s_net: std_logic_vector(25 downto 0);
  signal din: std_logic_vector(25 downto 0);
  signal dividend_data: std_logic_vector(25 downto 0);
  signal dividend_ready: std_logic;
  signal dividend_ready_x0: std_logic;
  signal dividend_valid_x0: std_logic;
  signal dividend_valid_x1: std_logic;
  signal dividend_valid_x2: std_logic;
  signal divider_dout_fracc: std_logic_vector(24 downto 0);
  signal divider_dout_valid_x0: std_logic;
  signal divisor_data: std_logic_vector(25 downto 0);
  signal divisor_data_x0: std_logic_vector(25 downto 0);
  signal divisor_ready: std_logic;
  signal divisor_valid_x0: std_logic;
  signal dout_down_x1: std_logic_vector(24 downto 0);
  signal dout_stretch: std_logic_vector(24 downto 0);
  signal down_sample1_q_net: std_logic_vector(24 downto 0);
  signal down_sample1_q_net_x26: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x27: std_logic_vector(23 downto 0);
  signal down_sample2_q_net: std_logic;
  signal down_sample2_q_net_x26: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x27: std_logic_vector(23 downto 0);
  signal down_sample3_q_net: std_logic_vector(24 downto 0);
  signal down_sample4_q_net: std_logic;
  signal down_sample5_q_net: std_logic_vector(24 downto 0);
  signal down_sample6_q_net: std_logic;
  signal down_sample7_q_net: std_logic_vector(24 downto 0);
  signal down_sample8_q_net: std_logic;
  signal down_sample_q_net: std_logic_vector(25 downto 0);
  signal expression1_dout_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical3_y_net_x2: std_logic;
  signal logical3_y_net_x3: std_logic;
  signal logical3_y_net_x4: std_logic;
  signal logical3_y_net_x5: std_logic;
  signal logical3_y_net_x6: std_logic;
  signal logical3_y_net_x7: std_logic;
  signal q_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal q_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal q_divider_s_axis_dividend_tready_net: std_logic;
  signal q_divider_s_axis_divisor_tready_net: std_logic;
  signal re_x0: std_logic;
  signal re_x1: std_logic;
  signal register10_q_net: std_logic_vector(25 downto 0);
  signal register11_q_net: std_logic_vector(24 downto 0);
  signal register12_q_net: std_logic_vector(24 downto 0);
  signal register13_q_net: std_logic_vector(24 downto 0);
  signal register14_q_net: std_logic_vector(25 downto 0);
  signal register1_q_net: std_logic_vector(24 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register1_q_net_x2: std_logic;
  signal register1_q_net_x3: std_logic;
  signal register1_q_net_x4: std_logic;
  signal register2_q_net: std_logic_vector(24 downto 0);
  signal register3_q_net: std_logic_vector(24 downto 0);
  signal register4_q_net: std_logic_vector(24 downto 0);
  signal register5_q_net: std_logic_vector(24 downto 0);
  signal register6_q_net: std_logic_vector(24 downto 0);
  signal register7_q_net: std_logic_vector(25 downto 0);
  signal register_q_net_x0: std_logic_vector(24 downto 0);
  signal register_q_net_x1: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(24 downto 0);
  signal register_q_net_x3: std_logic_vector(24 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret7_output_port_net: std_logic_vector(25 downto 0);
  signal reinterpret8_output_port_net: std_logic_vector(25 downto 0);
  signal relational_op_net: std_logic;
  signal sum_s_net: std_logic_vector(25 downto 0);
  signal up_sample2_q_net: std_logic_vector(25 downto 0);
  signal up_sample4_q_net: std_logic_vector(25 downto 0);
  signal up_sample6_q_net: std_logic_vector(25 downto 0);
  signal up_sample_q_net: std_logic_vector(25 downto 0);
  signal valid_ds_down_x1: std_logic;
  signal x_divider_m_axis_dout_tdata_fractional_net: std_logic_vector(24 downto 0);
  signal x_divider_m_axis_dout_tvalid_net_x0: std_logic;
  signal x_divider_s_axis_divisor_tready_net: std_logic;

begin
  down_sample2_q_net_x26 <= a;
  down_sample1_q_net_x26 <= b;
  down_sample2_q_net_x27 <= c;
  ce_1_sg_x90 <= ce_1;
  ce_2_sg_x37 <= ce_2;
  ce_70_sg_x26 <= ce_70;
  ce_logic_70_sg_x0 <= ce_logic_70;
  clk_1_sg_x90 <= clk_1;
  clk_2_sg_x37 <= clk_2;
  clk_70_sg_x26 <= clk_70;
  down_sample1_q_net_x27 <= d;
  del_sig_div_tbt_thres_i_net_x0 <= ds_thres;
  q <= assert8_dout_net_x1;
  q_valid <= assert9_dout_net_x1;
  sum_valid <= assert12_dout_net_x1;
  sum_x0 <= assert11_dout_net_x1;
  x <= assert5_dout_net_x1;
  x_valid <= assert10_dout_net_x1;
  y <= dout_down_x1;
  y_valid <= valid_ds_down_x1;

  a_plus_b: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x26,
      b => down_sample1_q_net_x26,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => a_plus_b_s_net
    );

  a_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x26,
      b => down_sample2_q_net_x27,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => a_plus_c_s_net
    );

  a_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x26,
      b => down_sample1_q_net_x27,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => a_plus_d_s_net
    );

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => q_divider_s_axis_dividend_tready_net,
      dout(0) => assert1_dout_net_x0
    );

  assert10: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample6_q_net,
      dout(0) => assert10_dout_net_x1
    );

  assert11: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample7_q_net,
      dout => assert11_dout_net_x1
    );

  assert12: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample8_q_net,
      dout(0) => assert12_dout_net_x1
    );

  assert2: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready_x0,
      dout(0) => re_x0
    );

  assert3: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => dividend_ready,
      dout(0) => re_x1
    );

  assert4: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample1_q_net,
      dout => dout_down_x1
    );

  assert5: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample5_q_net,
      dout => assert5_dout_net_x1
    );

  assert6: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => expression1_dout_net,
      dout(0) => assert6_dout_net_x0
    );

  assert7: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample2_q_net,
      dout(0) => valid_ds_down_x1
    );

  assert8: entity work.xlpassthrough
    generic map (
      din_width => 25,
      dout_width => 25
    )
    port map (
      din => down_sample3_q_net,
      dout => assert8_dout_net_x1
    );

  assert9: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => down_sample4_q_net,
      dout(0) => assert9_dout_net_x1
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => relational_op_net,
      dout(0) => assert_dout_net
    );

  b_plus_c: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x26,
      b => down_sample2_q_net_x27,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => b_plus_c_s_net
    );

  b_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample1_q_net_x26,
      b => down_sample1_q_net_x27,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => b_plus_d_s_net
    );

  c_plus_d: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 24,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 24,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 25,
      core_name0 => "addsb_11_0_293aa5f110d040c2",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 25,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 25
    )
    port map (
      a => down_sample2_q_net_x27,
      b => down_sample1_q_net_x27,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => c_plus_d_s_net
    );

  ce1: entity work.xlceprobe
    generic map (
      d_width => 1,
      q_width => 1
    )
    port map (
      ce => ce_logic_70_sg_x0,
      clk => clk_70_sg_x26,
      d(0) => assert_dout_net,
      q(0) => ce_70_x3
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 22,
      din_width => 26,
      dout_arith => 2,
      dout_bin_pt => 21,
      dout_width => 25,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlRound
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      clr => '0',
      din => delay_q_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  datareg_en1_e5d0399944: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      din => reinterpret2_output_port_net_x0,
      en => q_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x1,
      valid => register1_q_net_x2
    );

  datareg_en2_02a2053e69: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      din => reinterpret3_output_port_net_x0,
      en => x_divider_m_axis_dout_tvalid_net_x0,
      dout => register_q_net_x2,
      valid => register1_q_net_x3
    );

  datareg_en3_78179f99cc: entity work.datareg_en3_entity_6643090018
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      din => convert_dout_net_x0,
      en => delay1_q_net_x0,
      dout => register_q_net_x3,
      valid => register1_q_net_x4
    );

  datareg_en_ed948c360a: entity work.datareg_en_entity_79473f9ed1
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      din => reinterpret1_output_port_net_x0,
      en => divider_dout_valid_x0,
      dout => register_q_net_x0,
      valid => register1_q_net_x1
    );

  delay: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 26
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d => reinterpret8_output_port_net,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 56,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d(0) => logical3_y_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  delta_q: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register5_q_net,
      b => register6_q_net,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => delta_q_s_net
    );

  delta_x: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register1_q_net,
      b => register3_q_net,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => delta_x_s_net
    );

  delta_y: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_44053abf11139d96",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register2_q_net,
      b => register4_q_net,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => delta_y_s_net
    );

  down_sample: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      ds_ratio => 35,
      latency => 1,
      phase => 34,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register14_q_net,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_2_sg_x37,
      src_clk => clk_2_sg_x37,
      src_clr => '0',
      q => down_sample_q_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => dout_stretch,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q => down_sample1_q_net
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x0,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q(0) => down_sample2_q_net
    );

  down_sample3: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => register11_q_net,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q => down_sample3_q_net
    );

  down_sample4: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x1,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q(0) => down_sample4_q_net
    );

  down_sample5: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 24,
      d_width => 25,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlSigned,
      q_bin_pt => 24,
      q_width => 25
    )
    port map (
      d => register12_q_net,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q => down_sample5_q_net
    );

  down_sample6: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x2,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q(0) => down_sample6_q_net
    );

  down_sample7: entity work.xldsamp
    generic map (
      d_arith => xlSigned,
      d_bin_pt => 21,
      d_width => 25,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlSigned,
      q_bin_pt => 21,
      q_width => 25
    )
    port map (
      d => register13_q_net,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q => down_sample7_q_net
    );

  down_sample8: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      ds_ratio => 70,
      latency => 1,
      phase => 69,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => logical3_y_net_x3,
      dest_ce => ce_70_sg_x26,
      dest_clk => clk_70_sg_x26,
      dest_clr => '0',
      en => "1",
      src_ce => ce_1_sg_x90,
      src_clk => clk_1_sg_x90,
      src_clr => '0',
      q(0) => down_sample8_q_net
    );

  expression1: entity work.expr_375d7bbece
    port map (
      a(0) => x_divider_s_axis_divisor_tready_net,
      b(0) => divisor_ready,
      c(0) => q_divider_s_axis_divisor_tready_net,
      ce => '0',
      clk => '0',
      clr => '0',
      dout(0) => expression1_dout_net
    );

  pulse_stretcher1_eef5ee33be: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x2,
      extd_out => logical3_y_net_x1
    );

  pulse_stretcher2_6f5c3f41cf: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x3,
      extd_out => logical3_y_net_x2
    );

  pulse_stretcher3_e720dfd76f: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x4,
      extd_out => logical3_y_net_x3
    );

  pulse_stretcher4_0a5eb3f903: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => assert6_dout_net_x0,
      pulse_in => divisor_valid_x0,
      extd_out => logical3_y_net_x4
    );

  pulse_stretcher5_b95a604b09: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => re_x0,
      pulse_in => dividend_valid_x0,
      extd_out => logical3_y_net_x5
    );

  pulse_stretcher6_e7fb2961d9: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => assert1_dout_net_x0,
      pulse_in => dividend_valid_x1,
      extd_out => logical3_y_net_x6
    );

  pulse_stretcher7_6e7eb70147: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => re_x1,
      pulse_in => dividend_valid_x2,
      extd_out => logical3_y_net_x7
    );

  pulse_stretcher_f661707a58: entity work.pulse_stretcher_entity_9893378b63
    port map (
      ce_1 => ce_1_sg_x90,
      clk_1 => clk_1_sg_x90,
      clr => ce_70_x3,
      pulse_in => register1_q_net_x1,
      extd_out => logical3_y_net_x0
    );

  q_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      s_axis_dividend_tdata_dividend => reinterpret7_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x6,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => q_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => q_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => q_divider_s_axis_dividend_tready_net,
      s_axis_divisor_tready => q_divider_s_axis_divisor_tready_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => b_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register1_q_net
    );

  register10: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => delta_q_s_net,
      en => "1",
      rst => "0",
      q => register10_q_net
    );

  register11: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d => register_q_net_x1,
      en => "1",
      rst => "0",
      q => register11_q_net
    );

  register12: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d => register_q_net_x2,
      en => "1",
      rst => "0",
      q => register12_q_net
    );

  register13: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d => register_q_net_x3,
      en => "1",
      rst => "0",
      q => register13_q_net
    );

  register14: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_2_sg_x37,
      clk => clk_2_sg_x37,
      d => del_sig_div_tbt_thres_i_net_x0,
      en => "1",
      rst => "0",
      q => register14_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => a_plus_b_s_net,
      en => "1",
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => a_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => c_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => a_plus_c_s_net,
      en => "1",
      rst => "0",
      q => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => b_plus_d_s_net,
      en => "1",
      rst => "0",
      q => register6_q_net
    );

  register7: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => delta_x_s_net,
      en => "1",
      rst => "0",
      q => register7_q_net
    );

  register8: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => sum_s_net,
      en => "1",
      rst => "0",
      q => divisor_data
    );

  register9: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      d => delta_y_s_net,
      en => "1",
      rst => "0",
      q => din
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      d => register_q_net_x0,
      en => "1",
      rst => "0",
      q => dout_stretch
    );

  reinterpret1: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divider_dout_fracc,
      output_port => reinterpret1_output_port_net_x0
    );

  reinterpret2: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => q_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret2_output_port_net_x0
    );

  reinterpret3: entity work.reinterpret_31a4235b32
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => x_divider_m_axis_dout_tdata_fractional_net,
      output_port => reinterpret3_output_port_net_x0
    );

  reinterpret4: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample6_q_net,
      output_port => reinterpret4_output_port_net
    );

  reinterpret5: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample2_q_net,
      output_port => divisor_data_x0
    );

  reinterpret6: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample_q_net,
      output_port => dividend_data
    );

  reinterpret7: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => up_sample4_q_net,
      output_port => reinterpret7_output_port_net
    );

  reinterpret8: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => divisor_data_x0,
      output_port => reinterpret8_output_port_net
    );

  relational: entity work.relational_416cfcae1e
    port map (
      a => divisor_data,
      b => down_sample_q_net,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      op(0) => relational_op_net
    );

  sum: entity work.xladdsub
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 22,
      a_width => 25,
      b_arith => xlSigned,
      b_bin_pt => 22,
      b_width => 25,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 26,
      core_name0 => "addsb_11_0_3537d66a2361cd1e",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 26,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 22,
      s_width => 26
    )
    port map (
      a => register3_q_net,
      b => register1_q_net,
      ce => ce_70_sg_x26,
      clk => clk_70_sg_x26,
      clr => '0',
      en => "1",
      s => sum_s_net
    );

  up_sample: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => din,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q => up_sample_q_net
    );

  up_sample1: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q(0) => dividend_valid_x0
    );

  up_sample2: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => divisor_data,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q => up_sample2_q_net
    );

  up_sample3: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q(0) => divisor_valid_x0
    );

  up_sample4: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register10_q_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q => up_sample4_q_net
    );

  up_sample5: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q(0) => dividend_valid_x1
    );

  up_sample6: entity work.xlusamp
    generic map (
      copy_samples => 1,
      d_arith => xlSigned,
      d_bin_pt => 22,
      d_width => 26,
      latency => 0,
      q_arith => xlSigned,
      q_bin_pt => 22,
      q_width => 26
    )
    port map (
      d => register7_q_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q => up_sample6_q_net
    );

  up_sample7: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => assert_dout_net,
      dest_ce => ce_1_sg_x90,
      dest_clk => clk_1_sg_x90,
      dest_clr => '0',
      en => "1",
      src_ce => ce_70_sg_x26,
      src_clk => clk_70_sg_x26,
      src_clr => '0',
      q(0) => dividend_valid_x2
    );

  x_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      s_axis_dividend_tdata_dividend => reinterpret4_output_port_net,
      s_axis_dividend_tvalid => logical3_y_net_x7,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => x_divider_m_axis_dout_tdata_fractional_net,
      m_axis_dout_tvalid => x_divider_m_axis_dout_tvalid_net_x0,
      s_axis_dividend_tready => dividend_ready,
      s_axis_divisor_tready => x_divider_s_axis_divisor_tready_net
    );

  y_divider: entity work.xldivider_generator_47dc3a44bd8d9df86e42dac34ee6a9fc
    port map (
      ce => ce_1_sg_x90,
      clk => clk_1_sg_x90,
      s_axis_dividend_tdata_dividend => dividend_data,
      s_axis_dividend_tvalid => logical3_y_net_x5,
      s_axis_divisor_tdata_divisor => divisor_data_x0,
      s_axis_divisor_tvalid => logical3_y_net_x4,
      m_axis_dout_tdata_fractional => divider_dout_fracc,
      m_axis_dout_tvalid => divider_dout_valid_x0,
      s_axis_dividend_tready => dividend_ready_x0,
      s_axis_divisor_tready => divisor_ready
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/monit_pos_1/Cast1/format1"

entity format1_entity_a98b06306e is
  port (
    ce_56000000: in std_logic;
    clk_56000000: in std_logic;
    din: in std_logic_vector(25 downto 0);
    dout: out std_logic_vector(24 downto 0)
  );
end format1_entity_a98b06306e;

architecture structural of format1_entity_a98b06306e is
  signal ce_56000000_sg_x0: std_logic;
  signal clk_56000000_sg_x0: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal monit_pos_1_c_m_axis_data_tdata_net_x0: std_logic_vector(25 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(25 downto 0);

begin
  ce_56000000_sg_x0 <= ce_56000000;
  clk_56000000_sg_x0 <= clk_56000000;
  monit_pos_1_c_m_axis_data_tdata_net_x0 <= din;
  dout <= convert_dout_net_x0;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 24,
      din_width => 26,
      dout_arith => 2,
      dout_bin_pt => 24,
      dout_width => 25,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_56000000_sg_x0,
      clk => clk_56000000_sg_x0,
      clr => '0',
      din => reinterpret_output_port_net,
      en => "1",
      dout => convert_dout_net_x0
    );

  reinterpret: entity work.reinterpret_040ef1b598
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => monit_pos_1_c_m_axis_data_tdata_net_x0,
      output_port => reinterpret_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/monit_pos_1/Cast1"

entity cast1_entity_3d447d0833 is
  port (
    ce_56000000: in std_logic;
    clk_56000000: in std_logic;
    data_in: in std_logic_vector(25 downto 0);
    en: in std_logic;
    out_x0: out std_logic_vector(24 downto 0);
    vld_out: out std_logic
  );
end cast1_entity_3d447d0833;

architecture structural of cast1_entity_3d447d0833 is
  signal ce_56000000_sg_x1: std_logic;
  signal clk_56000000_sg_x1: std_logic;
  signal convert_dout_net_x0: std_logic_vector(24 downto 0);
  signal monit_pos_1_c_m_axis_data_tdata_net_x1: std_logic_vector(25 downto 0);
  signal monit_pos_1_c_m_axis_data_tvalid_net_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(24 downto 0);

begin
  ce_56000000_sg_x1 <= ce_56000000;
  clk_56000000_sg_x1 <= clk_56000000;
  monit_pos_1_c_m_axis_data_tdata_net_x1 <= data_in;
  monit_pos_1_c_m_axis_data_tvalid_net_x0 <= en;
  out_x0 <= register_q_net_x0;
  vld_out <= register1_q_net_x0;

  format1_a98b06306e: entity work.format1_entity_a98b06306e
    port map (
      ce_56000000 => ce_56000000_sg_x1,
      clk_56000000 => clk_56000000_sg_x1,
      din => monit_pos_1_c_m_axis_data_tdata_net_x1,
      dout => convert_dout_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_56000000_sg_x1,
      clk => clk_56000000_sg_x1,
      d(0) => monit_pos_1_c_m_axis_data_tvalid_net_x0,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 25,
      init_value => b"0000000000000000000000000"
    )
    port map (
      ce => ce_56000000_sg_x1,
      clk => clk_56000000_sg_x1,
      d => convert_dout_net_x0,
      en(0) => monit_pos_1_c_m_axis_data_tvalid_net_x0,
      rst => "0",
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/monit_pos_1/TDDM_monit_pos_1_out/TDDM_monit_pos_1_out_int"

entity tddm_monit_pos_1_out_int_entity_3405798202 is
  port (
    ce_224000000: in std_logic;
    ce_56000000: in std_logic;
    ch_in: in std_logic_vector(1 downto 0);
    clk_224000000: in std_logic;
    clk_56000000: in std_logic;
    din: in std_logic_vector(25 downto 0);
    dout_ch0: out std_logic_vector(25 downto 0);
    dout_ch1: out std_logic_vector(25 downto 0);
    dout_ch2: out std_logic_vector(25 downto 0);
    dout_ch3: out std_logic_vector(25 downto 0)
  );
end tddm_monit_pos_1_out_int_entity_3405798202;

architecture structural of tddm_monit_pos_1_out_int_entity_3405798202 is
  signal ce_224000000_sg_x4: std_logic;
  signal ce_56000000_sg_x2: std_logic;
  signal clk_224000000_sg_x4: std_logic;
  signal clk_56000000_sg_x2: std_logic;
  signal concat_y_net_x0: std_logic_vector(25 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal constant4_op_net: std_logic_vector(1 downto 0);
  signal constant_op_net: std_logic_vector(1 downto 0);
  signal down_sample1_q_net_x0: std_logic_vector(25 downto 0);
  signal down_sample2_q_net_x0: std_logic_vector(25 downto 0);
  signal down_sample3_q_net_x0: std_logic_vector(25 downto 0);
  signal down_sample4_q_net_x0: std_logic_vector(25 downto 0);
  signal register1_q_net: std_logic_vector(25 downto 0);
  signal register2_q_net: std_logic_vector(25 downto 0);
  signal register3_q_net: std_logic_vector(25 downto 0);
  signal register_q_net_x0: std_logic_vector(25 downto 0);
  signal register_q_net_x1: std_logic_vector(1 downto 0);
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational_op_net: std_logic;

begin
  ce_224000000_sg_x4 <= ce_224000000;
  ce_56000000_sg_x2 <= ce_56000000;
  register_q_net_x1 <= ch_in;
  clk_224000000_sg_x4 <= clk_224000000;
  clk_56000000_sg_x2 <= clk_56000000;
  concat_y_net_x0 <= din;
  dout_ch0 <= down_sample2_q_net_x0;
  dout_ch1 <= down_sample1_q_net_x0;
  dout_ch2 <= down_sample3_q_net_x0;
  dout_ch3 <= down_sample4_q_net_x0;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant3: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_e8ddc079e9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant_x0: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  down_sample1: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => register1_q_net,
      dest_ce => ce_224000000_sg_x4,
      dest_clk => clk_224000000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_56000000_sg_x2,
      src_clk => clk_56000000_sg_x2,
      src_clr => '0',
      q => down_sample1_q_net_x0
    );

  down_sample2: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => register_q_net_x0,
      dest_ce => ce_224000000_sg_x4,
      dest_clk => clk_224000000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_56000000_sg_x2,
      src_clk => clk_56000000_sg_x2,
      src_clr => '0',
      q => down_sample2_q_net_x0
    );

  down_sample3: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => register2_q_net,
      dest_ce => ce_224000000_sg_x4,
      dest_clk => clk_224000000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_56000000_sg_x2,
      src_clk => clk_56000000_sg_x2,
      src_clr => '0',
      q => down_sample3_q_net_x0
    );

  down_sample4: entity work.xldsamp
    generic map (
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 26,
      ds_ratio => 4,
      latency => 1,
      phase => 3,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 26
    )
    port map (
      d => register3_q_net,
      dest_ce => ce_224000000_sg_x4,
      dest_clk => clk_224000000_sg_x4,
      dest_clr => '0',
      en => "1",
      src_ce => ce_56000000_sg_x2,
      src_clk => clk_56000000_sg_x2,
      src_clr => '0',
      q => down_sample4_q_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      d => concat_y_net_x0,
      en(0) => relational1_op_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      d => concat_y_net_x0,
      en(0) => relational2_op_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      d => concat_y_net_x0,
      en(0) => relational3_op_net,
      rst => "0",
      q => register3_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 26,
      init_value => b"00000000000000000000000000"
    )
    port map (
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      d => concat_y_net_x0,
      en(0) => relational_op_net,
      rst => "0",
      q => register_q_net_x0
    );

  relational: entity work.relational_367321bc0c
    port map (
      a => register_q_net_x1,
      b => constant_op_net,
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_367321bc0c
    port map (
      a => register_q_net_x1,
      b => constant1_op_net,
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_367321bc0c
    port map (
      a => register_q_net_x1,
      b => constant3_op_net,
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_367321bc0c
    port map (
      a => register_q_net_x1,
      b => constant4_op_net,
      ce => ce_56000000_sg_x2,
      clk => clk_56000000_sg_x2,
      clr => '0',
      op(0) => relational3_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/monit_pos_1/TDDM_monit_pos_1_out"

entity tddm_monit_pos_1_out_entity_1d58a51dbf is
  port (
    ce_224000000: in std_logic;
    ce_56000000: in std_logic;
    clk_224000000: in std_logic;
    clk_56000000: in std_logic;
    monit_pos_1_ch_in: in std_logic_vector(1 downto 0);
    monit_pos_1_din: in std_logic_vector(25 downto 0);
    monit_pos_1_q_out: out std_logic_vector(25 downto 0);
    monit_pos_1_sum_out: out std_logic_vector(25 downto 0);
    monit_pos_1_x_out: out std_logic_vector(25 downto 0);
    monit_pos_1_y_out: out std_logic_vector(25 downto 0)
  );
end tddm_monit_pos_1_out_entity_1d58a51dbf;

architecture structural of tddm_monit_pos_1_out_entity_1d58a51dbf is
  signal ce_224000000_sg_x5: std_logic;
  signal ce_56000000_sg_x3: std_logic;
  signal clk_224000000_sg_x5: std_logic;
  signal clk_56000000_sg_x3: std_logic;
  signal concat_y_net_x1: std_logic_vector(25 downto 0);
  signal down_sample1_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample2_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample3_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample4_q_net_x1: std_logic_vector(25 downto 0);
  signal register_q_net_x2: std_logic_vector(1 downto 0);

begin
  ce_224000000_sg_x5 <= ce_224000000;
  ce_56000000_sg_x3 <= ce_56000000;
  clk_224000000_sg_x5 <= clk_224000000;
  clk_56000000_sg_x3 <= clk_56000000;
  register_q_net_x2 <= monit_pos_1_ch_in;
  concat_y_net_x1 <= monit_pos_1_din;
  monit_pos_1_q_out <= down_sample3_q_net_x1;
  monit_pos_1_sum_out <= down_sample4_q_net_x1;
  monit_pos_1_x_out <= down_sample2_q_net_x1;
  monit_pos_1_y_out <= down_sample1_q_net_x1;

  tddm_monit_pos_1_out_int_3405798202: entity work.tddm_monit_pos_1_out_int_entity_3405798202
    port map (
      ce_224000000 => ce_224000000_sg_x5,
      ce_56000000 => ce_56000000_sg_x3,
      ch_in => register_q_net_x2,
      clk_224000000 => clk_224000000_sg_x5,
      clk_56000000 => clk_56000000_sg_x3,
      din => concat_y_net_x1,
      dout_ch0 => down_sample2_q_net_x1,
      dout_ch1 => down_sample1_q_net_x1,
      dout_ch2 => down_sample3_q_net_x1,
      dout_ch3 => down_sample4_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066/monit_pos_1"

entity monit_pos_1_entity_522c8cf08d is
  port (
    ce_1: in std_logic;
    ce_224000000: in std_logic;
    ce_5600000: in std_logic;
    ce_56000000: in std_logic;
    ce_logic_5600000: in std_logic;
    ch_in: in std_logic_vector(1 downto 0);
    clk_1: in std_logic;
    clk_224000000: in std_logic;
    clk_5600000: in std_logic;
    clk_56000000: in std_logic;
    din: in std_logic_vector(24 downto 0);
    monit_1_pos_q: out std_logic_vector(24 downto 0);
    monit_1_pos_x: out std_logic_vector(24 downto 0);
    monit_1_pos_y: out std_logic_vector(24 downto 0);
    monit_1_sum: out std_logic_vector(24 downto 0);
    monit_1_vld_q: out std_logic;
    monit_1_vld_sum: out std_logic;
    monit_1_vld_x: out std_logic;
    monit_1_vld_y: out std_logic;
    monit_pos_1_c_x0: out std_logic
  );
end monit_pos_1_entity_522c8cf08d;

architecture structural of monit_pos_1_entity_522c8cf08d is
  signal ce_1_sg_x91: std_logic;
  signal ce_224000000_sg_x6: std_logic;
  signal ce_56000000_sg_x4: std_logic;
  signal ce_5600000_sg_x11: std_logic;
  signal ce_logic_5600000_sg_x1: std_logic;
  signal clk_1_sg_x91: std_logic;
  signal clk_224000000_sg_x6: std_logic;
  signal clk_56000000_sg_x4: std_logic;
  signal clk_5600000_sg_x11: std_logic;
  signal concat_y_net_x1: std_logic_vector(25 downto 0);
  signal down_sample1_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample2_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample3_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample4_q_net_x1: std_logic_vector(25 downto 0);
  signal down_sample_q_net_x3: std_logic_vector(1 downto 0);
  signal extractor1_dout_net: std_logic_vector(24 downto 0);
  signal extractor1_vld_out_net: std_logic;
  signal extractor2_dout_net: std_logic_vector(24 downto 0);
  signal extractor2_vld_out_net: std_logic;
  signal extractor3_dout_net: std_logic_vector(24 downto 0);
  signal extractor3_vld_out_net: std_logic;
  signal extractor4_dout_net: std_logic_vector(24 downto 0);
  signal extractor4_vld_out_net: std_logic;
  signal monit_pos_1_c_event_s_data_chanid_incorrect_net_x0: std_logic;
  signal monit_pos_1_c_m_axis_data_tdata_net_x1: std_logic_vector(25 downto 0);
  signal monit_pos_1_c_m_axis_data_tuser_chanid_net: std_logic_vector(1 downto 0);
  signal monit_pos_1_c_m_axis_data_tvalid_net_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register_q_net_x0: std_logic_vector(24 downto 0);
  signal register_q_net_x2: std_logic_vector(1 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret5_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret5_output_port_net_x1: std_logic_vector(24 downto 0);
  signal ufix_to_bool1_dout_net_x1: std_logic;
  signal ufix_to_bool2_dout_net_x1: std_logic;
  signal ufix_to_bool3_dout_net_x1: std_logic;
  signal ufix_to_bool_dout_net_x1: std_logic;

begin
  ce_1_sg_x91 <= ce_1;
  ce_224000000_sg_x6 <= ce_224000000;
  ce_5600000_sg_x11 <= ce_5600000;
  ce_56000000_sg_x4 <= ce_56000000;
  ce_logic_5600000_sg_x1 <= ce_logic_5600000;
  down_sample_q_net_x3 <= ch_in;
  clk_1_sg_x91 <= clk_1;
  clk_224000000_sg_x6 <= clk_224000000;
  clk_5600000_sg_x11 <= clk_5600000;
  clk_56000000_sg_x4 <= clk_56000000;
  reinterpret5_output_port_net_x1 <= din;
  monit_1_pos_q <= reinterpret2_output_port_net_x1;
  monit_1_pos_x <= reinterpret3_output_port_net_x1;
  monit_1_pos_y <= reinterpret1_output_port_net_x1;
  monit_1_sum <= reinterpret4_output_port_net_x1;
  monit_1_vld_q <= ufix_to_bool2_dout_net_x1;
  monit_1_vld_sum <= ufix_to_bool3_dout_net_x1;
  monit_1_vld_x <= ufix_to_bool_dout_net_x1;
  monit_1_vld_y <= ufix_to_bool1_dout_net_x1;
  monit_pos_1_c_x0 <= monit_pos_1_c_event_s_data_chanid_incorrect_net_x0;

  cast1_3d447d0833: entity work.cast1_entity_3d447d0833
    port map (
      ce_56000000 => ce_56000000_sg_x4,
      clk_56000000 => clk_56000000_sg_x4,
      data_in => monit_pos_1_c_m_axis_data_tdata_net_x1,
      en => monit_pos_1_c_m_axis_data_tvalid_net_x0,
      out_x0 => register_q_net_x0,
      vld_out => register1_q_net_x0
    );

  concat: entity work.concat_43e7f055fa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => register1_q_net_x0,
      in1 => reinterpret5_output_port_net,
      y => concat_y_net_x1
    );

  extractor1: entity work.bitbasher_a756ba0096
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      din => down_sample3_q_net_x1,
      dout => extractor1_dout_net,
      vld_out(0) => extractor1_vld_out_net
    );

  extractor2: entity work.bitbasher_a756ba0096
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      din => down_sample1_q_net_x1,
      dout => extractor2_dout_net,
      vld_out(0) => extractor2_vld_out_net
    );

  extractor3: entity work.bitbasher_a756ba0096
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      din => down_sample4_q_net_x1,
      dout => extractor3_dout_net,
      vld_out(0) => extractor3_vld_out_net
    );

  extractor4: entity work.bitbasher_a756ba0096
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      din => down_sample2_q_net_x1,
      dout => extractor4_dout_net,
      vld_out(0) => extractor4_vld_out_net
    );

  monit_pos_1_c: entity work.xlfir_compiler_eebfed0cb0075aa32aca169bb967f58b
    port map (
      ce => ce_1_sg_x91,
      ce_5600000 => ce_5600000_sg_x11,
      ce_56000000 => ce_56000000_sg_x4,
      ce_logic_5600000 => ce_logic_5600000_sg_x1,
      clk => clk_1_sg_x91,
      clk_5600000 => clk_5600000_sg_x11,
      clk_56000000 => clk_56000000_sg_x4,
      clk_logic_5600000 => clk_5600000_sg_x11,
      s_axis_data_tdata => reinterpret5_output_port_net_x1,
      s_axis_data_tuser_chanid => down_sample_q_net_x3,
      src_ce => ce_5600000_sg_x11,
      src_clk => clk_5600000_sg_x11,
      event_s_data_chanid_incorrect => monit_pos_1_c_event_s_data_chanid_incorrect_net_x0,
      m_axis_data_tdata => monit_pos_1_c_m_axis_data_tdata_net_x1,
      m_axis_data_tuser_chanid => monit_pos_1_c_m_axis_data_tuser_chanid_net,
      m_axis_data_tvalid => monit_pos_1_c_m_axis_data_tvalid_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 2,
      init_value => b"00"
    )
    port map (
      ce => ce_56000000_sg_x4,
      clk => clk_56000000_sg_x4,
      d => monit_pos_1_c_m_axis_data_tuser_chanid_net,
      en => "1",
      rst => "0",
      q => register_q_net_x2
    );

  reinterpret1: entity work.reinterpret_60ea556961
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => extractor2_dout_net,
      output_port => reinterpret1_output_port_net_x1
    );

  reinterpret2: entity work.reinterpret_60ea556961
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => extractor1_dout_net,
      output_port => reinterpret2_output_port_net_x1
    );

  reinterpret3: entity work.reinterpret_60ea556961
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => extractor4_dout_net,
      output_port => reinterpret3_output_port_net_x1
    );

  reinterpret4: entity work.reinterpret_60ea556961
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => extractor3_dout_net,
      output_port => reinterpret4_output_port_net_x1
    );

  reinterpret5: entity work.reinterpret_c3c0e847be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => register_q_net_x0,
      output_port => reinterpret5_output_port_net
    );

  tddm_monit_pos_1_out_1d58a51dbf: entity work.tddm_monit_pos_1_out_entity_1d58a51dbf
    port map (
      ce_224000000 => ce_224000000_sg_x6,
      ce_56000000 => ce_56000000_sg_x4,
      clk_224000000 => clk_224000000_sg_x6,
      clk_56000000 => clk_56000000_sg_x4,
      monit_pos_1_ch_in => register_q_net_x2,
      monit_pos_1_din => concat_y_net_x1,
      monit_pos_1_q_out => down_sample3_q_net_x1,
      monit_pos_1_sum_out => down_sample4_q_net_x1,
      monit_pos_1_x_out => down_sample2_q_net_x1,
      monit_pos_1_y_out => down_sample1_q_net_x1
    );

  ufix_to_bool: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_224000000_sg_x6,
      clk => clk_224000000_sg_x6,
      clr => '0',
      din(0) => extractor4_vld_out_net,
      en => "1",
      dout(0) => ufix_to_bool_dout_net_x1
    );

  ufix_to_bool1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_224000000_sg_x6,
      clk => clk_224000000_sg_x6,
      clr => '0',
      din(0) => extractor2_vld_out_net,
      en => "1",
      dout(0) => ufix_to_bool1_dout_net_x1
    );

  ufix_to_bool2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_224000000_sg_x6,
      clk => clk_224000000_sg_x6,
      clr => '0',
      din(0) => extractor1_vld_out_net,
      en => "1",
      dout(0) => ufix_to_bool2_dout_net_x1
    );

  ufix_to_bool3: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlRound
    )
    port map (
      ce => ce_224000000_sg_x6,
      clk => clk_224000000_sg_x6,
      clr => '0',
      din(0) => extractor3_vld_out_net,
      en => "1",
      dout(0) => ufix_to_bool3_dout_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "ddc_bpm_476_066"

entity ddc_bpm_476_066 is
  port (
    adc_ch0_i: in std_logic_vector(15 downto 0);
    adc_ch1_i: in std_logic_vector(15 downto 0);
    adc_ch2_i: in std_logic_vector(15 downto 0);
    adc_ch3_i: in std_logic_vector(15 downto 0);
    ce_1: in std_logic;
    ce_10000: in std_logic;
    ce_1120: in std_logic;
    ce_1400000: in std_logic;
    ce_2: in std_logic;
    ce_2240: in std_logic;
    ce_22400000: in std_logic;
    ce_224000000: in std_logic;
    ce_2500: in std_logic;
    ce_2800000: in std_logic;
    ce_35: in std_logic;
    ce_4480: in std_logic;
    ce_44800000: in std_logic;
    ce_5000: in std_logic;
    ce_560: in std_logic;
    ce_5600000: in std_logic;
    ce_56000000: in std_logic;
    ce_70: in std_logic;
    ce_logic_1: in std_logic;
    ce_logic_1400000: in std_logic;
    ce_logic_2240: in std_logic;
    ce_logic_22400000: in std_logic;
    ce_logic_2800000: in std_logic;
    ce_logic_560: in std_logic;
    ce_logic_5600000: in std_logic;
    ce_logic_70: in std_logic;
    clk_1: in std_logic;
    clk_10000: in std_logic;
    clk_1120: in std_logic;
    clk_1400000: in std_logic;
    clk_2: in std_logic;
    clk_2240: in std_logic;
    clk_22400000: in std_logic;
    clk_224000000: in std_logic;
    clk_2500: in std_logic;
    clk_2800000: in std_logic;
    clk_35: in std_logic;
    clk_4480: in std_logic;
    clk_44800000: in std_logic;
    clk_5000: in std_logic;
    clk_560: in std_logic;
    clk_5600000: in std_logic;
    clk_56000000: in std_logic;
    clk_70: in std_logic;
    dds_config_valid_ch0_i: in std_logic;
    dds_config_valid_ch1_i: in std_logic;
    dds_config_valid_ch2_i: in std_logic;
    dds_config_valid_ch3_i: in std_logic;
    dds_pinc_ch0_i: in std_logic_vector(29 downto 0);
    dds_pinc_ch1_i: in std_logic_vector(29 downto 0);
    dds_pinc_ch2_i: in std_logic_vector(29 downto 0);
    dds_pinc_ch3_i: in std_logic_vector(29 downto 0);
    dds_poff_ch0_i: in std_logic_vector(29 downto 0);
    dds_poff_ch1_i: in std_logic_vector(29 downto 0);
    dds_poff_ch2_i: in std_logic_vector(29 downto 0);
    dds_poff_ch3_i: in std_logic_vector(29 downto 0);
    del_sig_div_fofb_thres_i: in std_logic_vector(25 downto 0);
    del_sig_div_monit_thres_i: in std_logic_vector(25 downto 0);
    del_sig_div_tbt_thres_i: in std_logic_vector(25 downto 0);
    ksum_i: in std_logic_vector(24 downto 0);
    kx_i: in std_logic_vector(24 downto 0);
    ky_i: in std_logic_vector(24 downto 0);
    adc_ch0_dbg_data_o: out std_logic_vector(15 downto 0);
    adc_ch1_dbg_data_o: out std_logic_vector(15 downto 0);
    adc_ch2_dbg_data_o: out std_logic_vector(15 downto 0);
    adc_ch3_dbg_data_o: out std_logic_vector(15 downto 0);
    bpf_ch0_o: out std_logic_vector(23 downto 0);
    bpf_ch1_o: out std_logic_vector(23 downto 0);
    bpf_ch2_o: out std_logic_vector(23 downto 0);
    bpf_ch3_o: out std_logic_vector(23 downto 0);
    cic_fofb_q_01_missing_o: out std_logic;
    cic_fofb_q_23_missing_o: out std_logic;
    fofb_amp_ch0_o: out std_logic_vector(23 downto 0);
    fofb_amp_ch1_o: out std_logic_vector(23 downto 0);
    fofb_amp_ch2_o: out std_logic_vector(23 downto 0);
    fofb_amp_ch3_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch0_i_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch0_q_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch1_i_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch1_q_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch2_i_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch2_q_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch3_i_o: out std_logic_vector(23 downto 0);
    fofb_decim_ch3_q_o: out std_logic_vector(23 downto 0);
    fofb_pha_ch0_o: out std_logic_vector(23 downto 0);
    fofb_pha_ch1_o: out std_logic_vector(23 downto 0);
    fofb_pha_ch2_o: out std_logic_vector(23 downto 0);
    fofb_pha_ch3_o: out std_logic_vector(23 downto 0);
    mix_ch0_i_o: out std_logic_vector(23 downto 0);
    mix_ch0_q_o: out std_logic_vector(23 downto 0);
    mix_ch1_i_o: out std_logic_vector(23 downto 0);
    mix_ch1_q_o: out std_logic_vector(23 downto 0);
    mix_ch2_i_o: out std_logic_vector(23 downto 0);
    mix_ch2_q_o: out std_logic_vector(23 downto 0);
    mix_ch3_i_o: out std_logic_vector(23 downto 0);
    mix_ch3_q_o: out std_logic_vector(23 downto 0);
    monit_amp_ch0_o: out std_logic_vector(23 downto 0);
    monit_amp_ch1_o: out std_logic_vector(23 downto 0);
    monit_amp_ch2_o: out std_logic_vector(23 downto 0);
    monit_amp_ch3_o: out std_logic_vector(23 downto 0);
    monit_cfir_incorrect_o: out std_logic;
    monit_cic_unexpected_o: out std_logic;
    monit_pfir_incorrect_o: out std_logic;
    monit_pos_1_incorrect_o: out std_logic;
    q_fofb_o: out std_logic_vector(25 downto 0);
    q_fofb_valid_o: out std_logic;
    q_monit_1_o: out std_logic_vector(25 downto 0);
    q_monit_1_valid_o: out std_logic;
    q_monit_o: out std_logic_vector(25 downto 0);
    q_monit_valid_o: out std_logic;
    q_tbt_o: out std_logic_vector(25 downto 0);
    q_tbt_valid_o: out std_logic;
    sum_fofb_o: out std_logic_vector(25 downto 0);
    sum_fofb_valid_o: out std_logic;
    sum_monit_1_o: out std_logic_vector(25 downto 0);
    sum_monit_1_valid_o: out std_logic;
    sum_monit_o: out std_logic_vector(25 downto 0);
    sum_monit_valid_o: out std_logic;
    sum_tbt_o: out std_logic_vector(25 downto 0);
    sum_tbt_valid_o: out std_logic;
    tbt_amp_ch0_o: out std_logic_vector(23 downto 0);
    tbt_amp_ch1_o: out std_logic_vector(23 downto 0);
    tbt_amp_ch2_o: out std_logic_vector(23 downto 0);
    tbt_amp_ch3_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch01_incorrect_o: out std_logic;
    tbt_decim_ch0_i_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch0_q_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch1_i_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch1_q_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch23_incorrect_o: out std_logic;
    tbt_decim_ch2_i_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch2_q_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch3_i_o: out std_logic_vector(23 downto 0);
    tbt_decim_ch3_q_o: out std_logic_vector(23 downto 0);
    tbt_pha_ch0_o: out std_logic_vector(23 downto 0);
    tbt_pha_ch1_o: out std_logic_vector(23 downto 0);
    tbt_pha_ch2_o: out std_logic_vector(23 downto 0);
    tbt_pha_ch3_o: out std_logic_vector(23 downto 0);
    x_fofb_o: out std_logic_vector(25 downto 0);
    x_fofb_valid_o: out std_logic;
    x_monit_1_o: out std_logic_vector(25 downto 0);
    x_monit_1_valid_o: out std_logic;
    x_monit_o: out std_logic_vector(25 downto 0);
    x_monit_valid_o: out std_logic;
    x_tbt_o: out std_logic_vector(25 downto 0);
    x_tbt_valid_o: out std_logic;
    y_fofb_o: out std_logic_vector(25 downto 0);
    y_fofb_valid_o: out std_logic;
    y_monit_1_o: out std_logic_vector(25 downto 0);
    y_monit_1_valid_o: out std_logic;
    y_monit_o: out std_logic_vector(25 downto 0);
    y_monit_valid_o: out std_logic;
    y_tbt_o: out std_logic_vector(25 downto 0);
    y_tbt_valid_o: out std_logic
  );
end ddc_bpm_476_066;

architecture structural of ddc_bpm_476_066 is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "ddc_bpm_476_066,sysgen_core,{clock_period=4.44116092,clocking=Clock_Enables,compilation=HDL_Netlist,sample_periods=1.00000000000 2.00000000000 35.00000000000 70.00000000000 560.00000000000 1120.00000000000 2240.00000000000 2500.00000000000 4480.00000000000 5000.00000000000 10000.00000000000 1400000.00000000000 2800000.00000000000 5600000.00000000000 22400000.00000000000 44800000.00000000000 56000000.00000000000 224000000.00000000000,testbench=0,total_blocks=3299,xilinx_adder_subtracter_block=30,xilinx_arithmetic_relational_operator_block=66,xilinx_assert_block=39,xilinx_bit_slice_extractor_block=20,xilinx_bitbasher_block=5,xilinx_bitwise_expression_evaluator_block=3,xilinx_black_box_block=1,xilinx_bus_concatenator_block=9,xilinx_bus_multiplexer_block=8,xilinx_cic_compiler_3_0_block=5,xilinx_clock_enable_probe_block=11,xilinx_complex_multiplier_5_0__block=2,xilinx_constant_block_block=83,xilinx_cordic_5_0_block=4,xilinx_counter_block=8,xilinx_delay_block=59,xilinx_divider_generator_4_0_block=9,xilinx_down_sampler_block=102,xilinx_fir_compiler_6_3_block=5,xilinx_gateway_in_block=22,xilinx_gateway_out_block=233,xilinx_inverter_block=24,xilinx_logical_block_block=72,xilinx_multiplier_block=16,xilinx_register_block=264,xilinx_sample_time_block_block=88,xilinx_system_generator_block=1,xilinx_type_converter_block=23,xilinx_type_reinterpreter_block=94,xilinx_up_sampler_block=52,xilinx_wavescope_block=2,}";

  signal adc_ch0_dbg_data_o_net: std_logic_vector(15 downto 0);
  signal adc_ch0_i_net: std_logic_vector(15 downto 0);
  signal adc_ch1_dbg_data_o_net: std_logic_vector(15 downto 0);
  signal adc_ch1_i_net: std_logic_vector(15 downto 0);
  signal adc_ch2_dbg_data_o_net: std_logic_vector(15 downto 0);
  signal adc_ch2_i_net: std_logic_vector(15 downto 0);
  signal adc_ch3_dbg_data_o_net: std_logic_vector(15 downto 0);
  signal adc_ch3_i_net: std_logic_vector(15 downto 0);
  signal assert10_dout_net_x1: std_logic;
  signal assert10_dout_net_x2: std_logic;
  signal assert10_dout_net_x3: std_logic;
  signal assert11_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert11_dout_net_x2: std_logic_vector(24 downto 0);
  signal assert11_dout_net_x3: std_logic_vector(24 downto 0);
  signal assert12_dout_net_x1: std_logic;
  signal assert12_dout_net_x2: std_logic;
  signal assert12_dout_net_x3: std_logic;
  signal assert4_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert5_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert5_dout_net_x2: std_logic_vector(24 downto 0);
  signal assert5_dout_net_x3: std_logic_vector(24 downto 0);
  signal assert8_dout_net_x1: std_logic_vector(24 downto 0);
  signal assert8_dout_net_x2: std_logic_vector(24 downto 0);
  signal assert9_dout_net_x1: std_logic;
  signal assert9_dout_net_x2: std_logic;
  signal assert9_dout_net_x3: std_logic;
  signal bpf_ch0_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch1_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch2_o_net: std_logic_vector(23 downto 0);
  signal bpf_ch3_o_net: std_logic_vector(23 downto 0);
  signal ce_10000_sg_x2: std_logic;
  signal ce_1120_sg_x32: std_logic;
  signal ce_1400000_sg_x3: std_logic;
  signal ce_1_sg_x92: std_logic;
  signal ce_224000000_sg_x7: std_logic;
  signal ce_22400000_sg_x28: std_logic;
  signal ce_2240_sg_x28: std_logic;
  signal ce_2500_sg_x3: std_logic;
  signal ce_2800000_sg_x4: std_logic;
  signal ce_2_sg_x38: std_logic;
  signal ce_35_sg_x22: std_logic;
  signal ce_44800000_sg_x2: std_logic;
  signal ce_4480_sg_x9: std_logic;
  signal ce_5000_sg_x9: std_logic;
  signal ce_56000000_sg_x5: std_logic;
  signal ce_5600000_sg_x12: std_logic;
  signal ce_560_sg_x3: std_logic;
  signal ce_70_sg_x27: std_logic;
  signal ce_logic_1400000_sg_x2: std_logic;
  signal ce_logic_1_sg_x20: std_logic;
  signal ce_logic_22400000_sg_x1: std_logic;
  signal ce_logic_2240_sg_x1: std_logic;
  signal ce_logic_2800000_sg_x2: std_logic;
  signal ce_logic_5600000_sg_x2: std_logic;
  signal ce_logic_560_sg_x3: std_logic;
  signal ce_logic_70_sg_x1: std_logic;
  signal ch_out_x2: std_logic_vector(1 downto 0);
  signal cic_fofb_q_01_missing_o_net: std_logic;
  signal cic_fofb_q_23_missing_o_net: std_logic;
  signal clk_10000_sg_x2: std_logic;
  signal clk_1120_sg_x32: std_logic;
  signal clk_1400000_sg_x3: std_logic;
  signal clk_1_sg_x92: std_logic;
  signal clk_224000000_sg_x7: std_logic;
  signal clk_22400000_sg_x28: std_logic;
  signal clk_2240_sg_x28: std_logic;
  signal clk_2500_sg_x3: std_logic;
  signal clk_2800000_sg_x4: std_logic;
  signal clk_2_sg_x38: std_logic;
  signal clk_35_sg_x22: std_logic;
  signal clk_44800000_sg_x2: std_logic;
  signal clk_4480_sg_x9: std_logic;
  signal clk_5000_sg_x9: std_logic;
  signal clk_56000000_sg_x5: std_logic;
  signal clk_5600000_sg_x12: std_logic;
  signal clk_560_sg_x3: std_logic;
  signal clk_70_sg_x27: std_logic;
  signal concat1_y_net_x0: std_logic_vector(25 downto 0);
  signal concat2_y_net_x0: std_logic_vector(25 downto 0);
  signal concat3_y_net_x0: std_logic_vector(25 downto 0);
  signal concat_y_net_x0: std_logic_vector(25 downto 0);
  signal constant10_op_net_x0: std_logic;
  signal constant11_op_net_x0: std_logic;
  signal constant15_op_net_x1: std_logic;
  signal constant3_op_net_x1: std_logic;
  signal dds_config_valid_ch0_i_net: std_logic;
  signal dds_config_valid_ch1_i_net: std_logic;
  signal dds_config_valid_ch2_i_net: std_logic;
  signal dds_config_valid_ch3_i_net: std_logic;
  signal dds_pinc_ch0_i_net: std_logic_vector(29 downto 0);
  signal dds_pinc_ch1_i_net: std_logic_vector(29 downto 0);
  signal dds_pinc_ch2_i_net: std_logic_vector(29 downto 0);
  signal dds_pinc_ch3_i_net: std_logic_vector(29 downto 0);
  signal dds_poff_ch0_i_net: std_logic_vector(29 downto 0);
  signal dds_poff_ch1_i_net: std_logic_vector(29 downto 0);
  signal dds_poff_ch2_i_net: std_logic_vector(29 downto 0);
  signal dds_poff_ch3_i_net: std_logic_vector(29 downto 0);
  signal del_sig_div_fofb_thres_i_net: std_logic_vector(25 downto 0);
  signal del_sig_div_monit_thres_i_net: std_logic_vector(25 downto 0);
  signal del_sig_div_tbt_thres_i_net: std_logic_vector(25 downto 0);
  signal dout_down_x1: std_logic_vector(24 downto 0);
  signal dout_down_x2: std_logic_vector(24 downto 0);
  signal dout_down_x3: std_logic_vector(24 downto 0);
  signal dout_x2: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x34: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x35: std_logic_vector(23 downto 0);
  signal down_sample1_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x20: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x21: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x34: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x35: std_logic_vector(23 downto 0);
  signal down_sample2_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample3_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample4_q_net_x5: std_logic_vector(23 downto 0);
  signal down_sample_q_net_x3: std_logic_vector(1 downto 0);
  signal down_sample_q_net_x4: std_logic_vector(25 downto 0);
  signal fofb_amp_ch0_o_net: std_logic_vector(23 downto 0);
  signal fofb_amp_ch1_o_net: std_logic_vector(23 downto 0);
  signal fofb_amp_ch2_o_net: std_logic_vector(23 downto 0);
  signal fofb_amp_ch3_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch0_i_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch0_q_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch1_i_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch1_q_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch2_i_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch2_q_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch3_i_o_net: std_logic_vector(23 downto 0);
  signal fofb_decim_ch3_q_o_net: std_logic_vector(23 downto 0);
  signal fofb_pha_ch0_o_net: std_logic_vector(23 downto 0);
  signal fofb_pha_ch1_o_net: std_logic_vector(23 downto 0);
  signal fofb_pha_ch2_o_net: std_logic_vector(23 downto 0);
  signal fofb_pha_ch3_o_net: std_logic_vector(23 downto 0);
  signal ksum_i_net: std_logic_vector(24 downto 0);
  signal kx_i_net: std_logic_vector(24 downto 0);
  signal ky_i_net: std_logic_vector(24 downto 0);
  signal mix_ch0_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch0_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch1_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch1_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch2_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch2_q_o_net: std_logic_vector(23 downto 0);
  signal mix_ch3_i_o_net: std_logic_vector(23 downto 0);
  signal mix_ch3_q_o_net: std_logic_vector(23 downto 0);
  signal monit_amp_ch0_o_net: std_logic_vector(23 downto 0);
  signal monit_amp_ch1_o_net: std_logic_vector(23 downto 0);
  signal monit_amp_ch2_o_net: std_logic_vector(23 downto 0);
  signal monit_amp_ch3_o_net: std_logic_vector(23 downto 0);
  signal monit_cfir_incorrect_o_net: std_logic;
  signal monit_cic_unexpected_o_net: std_logic;
  signal monit_pfir_incorrect_o_net: std_logic;
  signal monit_pos_1_incorrect_o_net: std_logic;
  signal q_fofb_o_net: std_logic_vector(25 downto 0);
  signal q_fofb_valid_o_net: std_logic;
  signal q_monit_1_o_net: std_logic_vector(25 downto 0);
  signal q_monit_1_valid_o_net: std_logic;
  signal q_monit_o_net: std_logic_vector(25 downto 0);
  signal q_monit_valid_o_net: std_logic;
  signal q_tbt_o_net: std_logic_vector(25 downto 0);
  signal q_tbt_valid_o_net: std_logic;
  signal register1_q_net_x6: std_logic;
  signal register1_q_net_x7: std_logic;
  signal register3_q_net_x15: std_logic;
  signal register3_q_net_x16: std_logic;
  signal register4_q_net_x14: std_logic_vector(23 downto 0);
  signal register4_q_net_x15: std_logic_vector(23 downto 0);
  signal register5_q_net_x11: std_logic_vector(23 downto 0);
  signal register5_q_net_x15: std_logic_vector(23 downto 0);
  signal register_q_net_x12: std_logic_vector(23 downto 0);
  signal register_q_net_x13: std_logic_vector(23 downto 0);
  signal register_q_net_x14: std_logic_vector(23 downto 0);
  signal register_q_net_x15: std_logic_vector(23 downto 0);
  signal register_q_net_x31: std_logic_vector(23 downto 0);
  signal register_q_net_x32: std_logic_vector(23 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net: std_logic_vector(24 downto 0);
  signal reinterpret4_output_port_net_x1: std_logic_vector(24 downto 0);
  signal reinterpret5_output_port_net_x1: std_logic_vector(24 downto 0);
  signal sum_fofb_o_net: std_logic_vector(25 downto 0);
  signal sum_fofb_valid_o_net: std_logic;
  signal sum_monit_1_o_net: std_logic_vector(25 downto 0);
  signal sum_monit_1_valid_o_net: std_logic;
  signal sum_monit_o_net: std_logic_vector(25 downto 0);
  signal sum_monit_valid_o_net: std_logic;
  signal sum_tbt_o_net: std_logic_vector(25 downto 0);
  signal sum_tbt_valid_o_net: std_logic;
  signal tbt_amp_ch0_o_net: std_logic_vector(23 downto 0);
  signal tbt_amp_ch1_o_net: std_logic_vector(23 downto 0);
  signal tbt_amp_ch2_o_net: std_logic_vector(23 downto 0);
  signal tbt_amp_ch3_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch01_incorrect_o_net: std_logic;
  signal tbt_decim_ch0_i_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch0_q_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch1_i_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch1_q_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch23_incorrect_o_net: std_logic;
  signal tbt_decim_ch2_i_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch2_q_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch3_i_o_net: std_logic_vector(23 downto 0);
  signal tbt_decim_ch3_q_o_net: std_logic_vector(23 downto 0);
  signal tbt_pha_ch0_o_net: std_logic_vector(23 downto 0);
  signal tbt_pha_ch1_o_net: std_logic_vector(23 downto 0);
  signal tbt_pha_ch2_o_net: std_logic_vector(23 downto 0);
  signal tbt_pha_ch3_o_net: std_logic_vector(23 downto 0);
  signal ufix_to_bool1_dout_net_x1: std_logic;
  signal ufix_to_bool2_dout_net_x1: std_logic;
  signal ufix_to_bool3_dout_net_x1: std_logic;
  signal ufix_to_bool_dout_net_x1: std_logic;
  signal valid_ds_down_x1: std_logic;
  signal valid_ds_down_x2: std_logic;
  signal valid_ds_down_x3: std_logic;
  signal x_fofb_o_net: std_logic_vector(25 downto 0);
  signal x_fofb_valid_o_net: std_logic;
  signal x_monit_1_o_net: std_logic_vector(25 downto 0);
  signal x_monit_1_valid_o_net: std_logic;
  signal x_monit_o_net: std_logic_vector(25 downto 0);
  signal x_monit_valid_o_net: std_logic;
  signal x_tbt_o_net: std_logic_vector(25 downto 0);
  signal x_tbt_valid_o_net: std_logic;
  signal y_fofb_o_net: std_logic_vector(25 downto 0);
  signal y_fofb_valid_o_net: std_logic;
  signal y_monit_1_o_net: std_logic_vector(25 downto 0);
  signal y_monit_1_valid_o_net: std_logic;
  signal y_monit_o_net: std_logic_vector(25 downto 0);
  signal y_monit_valid_o_net: std_logic;
  signal y_tbt_o_net: std_logic_vector(25 downto 0);
  signal y_tbt_valid_o_net: std_logic;

begin
  adc_ch0_i_net <= adc_ch0_i;
  adc_ch1_i_net <= adc_ch1_i;
  adc_ch2_i_net <= adc_ch2_i;
  adc_ch3_i_net <= adc_ch3_i;
  ce_1_sg_x92 <= ce_1;
  ce_10000_sg_x2 <= ce_10000;
  ce_1120_sg_x32 <= ce_1120;
  ce_1400000_sg_x3 <= ce_1400000;
  ce_2_sg_x38 <= ce_2;
  ce_2240_sg_x28 <= ce_2240;
  ce_22400000_sg_x28 <= ce_22400000;
  ce_224000000_sg_x7 <= ce_224000000;
  ce_2500_sg_x3 <= ce_2500;
  ce_2800000_sg_x4 <= ce_2800000;
  ce_35_sg_x22 <= ce_35;
  ce_4480_sg_x9 <= ce_4480;
  ce_44800000_sg_x2 <= ce_44800000;
  ce_5000_sg_x9 <= ce_5000;
  ce_560_sg_x3 <= ce_560;
  ce_5600000_sg_x12 <= ce_5600000;
  ce_56000000_sg_x5 <= ce_56000000;
  ce_70_sg_x27 <= ce_70;
  ce_logic_1_sg_x20 <= ce_logic_1;
  ce_logic_1400000_sg_x2 <= ce_logic_1400000;
  ce_logic_2240_sg_x1 <= ce_logic_2240;
  ce_logic_22400000_sg_x1 <= ce_logic_22400000;
  ce_logic_2800000_sg_x2 <= ce_logic_2800000;
  ce_logic_560_sg_x3 <= ce_logic_560;
  ce_logic_5600000_sg_x2 <= ce_logic_5600000;
  ce_logic_70_sg_x1 <= ce_logic_70;
  clk_1_sg_x92 <= clk_1;
  clk_10000_sg_x2 <= clk_10000;
  clk_1120_sg_x32 <= clk_1120;
  clk_1400000_sg_x3 <= clk_1400000;
  clk_2_sg_x38 <= clk_2;
  clk_2240_sg_x28 <= clk_2240;
  clk_22400000_sg_x28 <= clk_22400000;
  clk_224000000_sg_x7 <= clk_224000000;
  clk_2500_sg_x3 <= clk_2500;
  clk_2800000_sg_x4 <= clk_2800000;
  clk_35_sg_x22 <= clk_35;
  clk_4480_sg_x9 <= clk_4480;
  clk_44800000_sg_x2 <= clk_44800000;
  clk_5000_sg_x9 <= clk_5000;
  clk_560_sg_x3 <= clk_560;
  clk_5600000_sg_x12 <= clk_5600000;
  clk_56000000_sg_x5 <= clk_56000000;
  clk_70_sg_x27 <= clk_70;
  dds_config_valid_ch0_i_net <= dds_config_valid_ch0_i;
  dds_config_valid_ch1_i_net <= dds_config_valid_ch1_i;
  dds_config_valid_ch2_i_net <= dds_config_valid_ch2_i;
  dds_config_valid_ch3_i_net <= dds_config_valid_ch3_i;
  dds_pinc_ch0_i_net <= dds_pinc_ch0_i;
  dds_pinc_ch1_i_net <= dds_pinc_ch1_i;
  dds_pinc_ch2_i_net <= dds_pinc_ch2_i;
  dds_pinc_ch3_i_net <= dds_pinc_ch3_i;
  dds_poff_ch0_i_net <= dds_poff_ch0_i;
  dds_poff_ch1_i_net <= dds_poff_ch1_i;
  dds_poff_ch2_i_net <= dds_poff_ch2_i;
  dds_poff_ch3_i_net <= dds_poff_ch3_i;
  del_sig_div_fofb_thres_i_net <= del_sig_div_fofb_thres_i;
  del_sig_div_monit_thres_i_net <= del_sig_div_monit_thres_i;
  del_sig_div_tbt_thres_i_net <= del_sig_div_tbt_thres_i;
  ksum_i_net <= ksum_i;
  kx_i_net <= kx_i;
  ky_i_net <= ky_i;
  adc_ch0_dbg_data_o <= adc_ch0_dbg_data_o_net;
  adc_ch1_dbg_data_o <= adc_ch1_dbg_data_o_net;
  adc_ch2_dbg_data_o <= adc_ch2_dbg_data_o_net;
  adc_ch3_dbg_data_o <= adc_ch3_dbg_data_o_net;
  bpf_ch0_o <= bpf_ch0_o_net;
  bpf_ch1_o <= bpf_ch1_o_net;
  bpf_ch2_o <= bpf_ch2_o_net;
  bpf_ch3_o <= bpf_ch3_o_net;
  cic_fofb_q_01_missing_o <= cic_fofb_q_01_missing_o_net;
  cic_fofb_q_23_missing_o <= cic_fofb_q_23_missing_o_net;
  fofb_amp_ch0_o <= fofb_amp_ch0_o_net;
  fofb_amp_ch1_o <= fofb_amp_ch1_o_net;
  fofb_amp_ch2_o <= fofb_amp_ch2_o_net;
  fofb_amp_ch3_o <= fofb_amp_ch3_o_net;
  fofb_decim_ch0_i_o <= fofb_decim_ch0_i_o_net;
  fofb_decim_ch0_q_o <= fofb_decim_ch0_q_o_net;
  fofb_decim_ch1_i_o <= fofb_decim_ch1_i_o_net;
  fofb_decim_ch1_q_o <= fofb_decim_ch1_q_o_net;
  fofb_decim_ch2_i_o <= fofb_decim_ch2_i_o_net;
  fofb_decim_ch2_q_o <= fofb_decim_ch2_q_o_net;
  fofb_decim_ch3_i_o <= fofb_decim_ch3_i_o_net;
  fofb_decim_ch3_q_o <= fofb_decim_ch3_q_o_net;
  fofb_pha_ch0_o <= fofb_pha_ch0_o_net;
  fofb_pha_ch1_o <= fofb_pha_ch1_o_net;
  fofb_pha_ch2_o <= fofb_pha_ch2_o_net;
  fofb_pha_ch3_o <= fofb_pha_ch3_o_net;
  mix_ch0_i_o <= mix_ch0_i_o_net;
  mix_ch0_q_o <= mix_ch0_q_o_net;
  mix_ch1_i_o <= mix_ch1_i_o_net;
  mix_ch1_q_o <= mix_ch1_q_o_net;
  mix_ch2_i_o <= mix_ch2_i_o_net;
  mix_ch2_q_o <= mix_ch2_q_o_net;
  mix_ch3_i_o <= mix_ch3_i_o_net;
  mix_ch3_q_o <= mix_ch3_q_o_net;
  monit_amp_ch0_o <= monit_amp_ch0_o_net;
  monit_amp_ch1_o <= monit_amp_ch1_o_net;
  monit_amp_ch2_o <= monit_amp_ch2_o_net;
  monit_amp_ch3_o <= monit_amp_ch3_o_net;
  monit_cfir_incorrect_o <= monit_cfir_incorrect_o_net;
  monit_cic_unexpected_o <= monit_cic_unexpected_o_net;
  monit_pfir_incorrect_o <= monit_pfir_incorrect_o_net;
  monit_pos_1_incorrect_o <= monit_pos_1_incorrect_o_net;
  q_fofb_o <= q_fofb_o_net;
  q_fofb_valid_o <= q_fofb_valid_o_net;
  q_monit_1_o <= q_monit_1_o_net;
  q_monit_1_valid_o <= q_monit_1_valid_o_net;
  q_monit_o <= q_monit_o_net;
  q_monit_valid_o <= q_monit_valid_o_net;
  q_tbt_o <= q_tbt_o_net;
  q_tbt_valid_o <= q_tbt_valid_o_net;
  sum_fofb_o <= sum_fofb_o_net;
  sum_fofb_valid_o <= sum_fofb_valid_o_net;
  sum_monit_1_o <= sum_monit_1_o_net;
  sum_monit_1_valid_o <= sum_monit_1_valid_o_net;
  sum_monit_o <= sum_monit_o_net;
  sum_monit_valid_o <= sum_monit_valid_o_net;
  sum_tbt_o <= sum_tbt_o_net;
  sum_tbt_valid_o <= sum_tbt_valid_o_net;
  tbt_amp_ch0_o <= tbt_amp_ch0_o_net;
  tbt_amp_ch1_o <= tbt_amp_ch1_o_net;
  tbt_amp_ch2_o <= tbt_amp_ch2_o_net;
  tbt_amp_ch3_o <= tbt_amp_ch3_o_net;
  tbt_decim_ch01_incorrect_o <= tbt_decim_ch01_incorrect_o_net;
  tbt_decim_ch0_i_o <= tbt_decim_ch0_i_o_net;
  tbt_decim_ch0_q_o <= tbt_decim_ch0_q_o_net;
  tbt_decim_ch1_i_o <= tbt_decim_ch1_i_o_net;
  tbt_decim_ch1_q_o <= tbt_decim_ch1_q_o_net;
  tbt_decim_ch23_incorrect_o <= tbt_decim_ch23_incorrect_o_net;
  tbt_decim_ch2_i_o <= tbt_decim_ch2_i_o_net;
  tbt_decim_ch2_q_o <= tbt_decim_ch2_q_o_net;
  tbt_decim_ch3_i_o <= tbt_decim_ch3_i_o_net;
  tbt_decim_ch3_q_o <= tbt_decim_ch3_q_o_net;
  tbt_pha_ch0_o <= tbt_pha_ch0_o_net;
  tbt_pha_ch1_o <= tbt_pha_ch1_o_net;
  tbt_pha_ch2_o <= tbt_pha_ch2_o_net;
  tbt_pha_ch3_o <= tbt_pha_ch3_o_net;
  x_fofb_o <= x_fofb_o_net;
  x_fofb_valid_o <= x_fofb_valid_o_net;
  x_monit_1_o <= x_monit_1_o_net;
  x_monit_1_valid_o <= x_monit_1_valid_o_net;
  x_monit_o <= x_monit_o_net;
  x_monit_valid_o <= x_monit_valid_o_net;
  x_tbt_o <= x_tbt_o_net;
  x_tbt_valid_o <= x_tbt_valid_o_net;
  y_fofb_o <= y_fofb_o_net;
  y_fofb_valid_o <= y_fofb_valid_o_net;
  y_monit_1_o <= y_monit_1_o_net;
  y_monit_1_valid_o <= y_monit_1_valid_o_net;
  y_monit_o <= y_monit_o_net;
  y_monit_valid_o <= y_monit_valid_o_net;
  y_tbt_o <= y_tbt_o_net;
  y_tbt_valid_o <= y_tbt_valid_o_net;

  bpf_d31c4af409: entity work.bpf_entity_d31c4af409
    port map (
      din_ch0 => adc_ch0_dbg_data_o_net,
      din_ch1 => adc_ch1_dbg_data_o_net,
      din_ch2 => adc_ch2_dbg_data_o_net,
      din_ch3 => adc_ch3_dbg_data_o_net,
      dout_ch0 => bpf_ch0_o_net,
      dout_ch1 => bpf_ch1_o_net,
      dout_ch2 => bpf_ch2_o_net,
      dout_ch3 => bpf_ch3_o_net
    );

  concat: entity work.concat_43e7f055fa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => assert12_dout_net_x2,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net_x0
    );

  concat1: entity work.concat_43e7f055fa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => valid_ds_down_x2,
      in1 => reinterpret2_output_port_net,
      y => concat1_y_net_x0
    );

  concat2: entity work.concat_43e7f055fa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => assert9_dout_net_x2,
      in1 => reinterpret3_output_port_net,
      y => concat2_y_net_x0
    );

  concat3: entity work.concat_43e7f055fa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => assert10_dout_net_x2,
      in1 => reinterpret4_output_port_net,
      y => concat3_y_net_x0
    );

  constant10: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant10_op_net_x0
    );

  constant11: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant11_op_net_x0
    );

  constant15: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant15_op_net_x1
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net_x1
    );

  convert_filt_fda412c1bf: entity work.convert_filt_entity_fda412c1bf
    port map (
      din => down_sample_q_net_x4,
      dout => reinterpret5_output_port_net_x1
    );

  dds_sub_a4b6b880f6: entity work.dds_sub_entity_a4b6b880f6
    port map (
      ce_1 => ce_1_sg_x92,
      ce_2 => ce_2_sg_x38,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x92,
      clk_2 => clk_2_sg_x38,
      dds_01_cosine => register_q_net_x12,
      dds_01_sine => register_q_net_x13,
      dds_23_cosine => register_q_net_x14,
      dds_23_sine => register_q_net_x15
    );

  delta_sigma_fofb_ee61e649ea: entity work.delta_sigma_fofb_entity_ee61e649ea
    port map (
      a => down_sample2_q_net_x20,
      b => down_sample1_q_net_x20,
      c => down_sample2_q_net_x21,
      ce_1 => ce_1_sg_x92,
      ce_2 => ce_2_sg_x38,
      ce_2240 => ce_2240_sg_x28,
      ce_logic_2240 => ce_logic_2240_sg_x1,
      clk_1 => clk_1_sg_x92,
      clk_2 => clk_2_sg_x38,
      clk_2240 => clk_2240_sg_x28,
      d => down_sample1_q_net_x21,
      ds_thres => del_sig_div_fofb_thres_i_net,
      q => assert8_dout_net_x1,
      q_valid => assert9_dout_net_x1,
      sum_valid => assert12_dout_net_x1,
      sum_x0 => assert11_dout_net_x1,
      x => assert5_dout_net_x1,
      x_valid => assert10_dout_net_x1,
      y => dout_down_x1,
      y_valid => valid_ds_down_x1
    );

  delta_sigma_monit_a8f8b81626: entity work.delta_sigma_monit_entity_a8f8b81626
    port map (
      a => down_sample2_q_net_x5,
      b => down_sample1_q_net_x5,
      c => down_sample3_q_net_x5,
      ce_1 => ce_1_sg_x92,
      ce_10000 => ce_10000_sg_x2,
      ce_2 => ce_2_sg_x38,
      ce_22400000 => ce_22400000_sg_x28,
      ce_4480 => ce_4480_sg_x9,
      ce_44800000 => ce_44800000_sg_x2,
      ce_5000 => ce_5000_sg_x9,
      ce_logic_22400000 => ce_logic_22400000_sg_x1,
      clk_1 => clk_1_sg_x92,
      clk_10000 => clk_10000_sg_x2,
      clk_2 => clk_2_sg_x38,
      clk_22400000 => clk_22400000_sg_x28,
      clk_4480 => clk_4480_sg_x9,
      clk_44800000 => clk_44800000_sg_x2,
      clk_5000 => clk_5000_sg_x9,
      d => down_sample4_q_net_x5,
      ds_thres => del_sig_div_monit_thres_i_net,
      q => assert4_dout_net_x1,
      q_valid => assert9_dout_net_x2,
      sum_valid => assert10_dout_net_x2,
      sum_x0 => assert5_dout_net_x2,
      x => assert11_dout_net_x2,
      x_valid => assert12_dout_net_x2,
      y => dout_down_x2,
      y_valid => valid_ds_down_x2
    );

  delta_sigma_tbt_bbfa8a8a69: entity work.delta_sigma_tbt_entity_bbfa8a8a69
    port map (
      a => down_sample2_q_net_x34,
      b => down_sample1_q_net_x34,
      c => down_sample2_q_net_x35,
      ce_1 => ce_1_sg_x92,
      ce_2 => ce_2_sg_x38,
      ce_70 => ce_70_sg_x27,
      ce_logic_70 => ce_logic_70_sg_x1,
      clk_1 => clk_1_sg_x92,
      clk_2 => clk_2_sg_x38,
      clk_70 => clk_70_sg_x27,
      d => down_sample1_q_net_x35,
      ds_thres => del_sig_div_tbt_thres_i_net,
      q => assert8_dout_net_x2,
      q_valid => assert9_dout_net_x3,
      sum_valid => assert12_dout_net_x3,
      sum_x0 => assert11_dout_net_x3,
      x => assert5_dout_net_x3,
      x_valid => assert10_dout_net_x3,
      y => dout_down_x3,
      y_valid => valid_ds_down_x3
    );

  fofb_amp_8b25d4b0b6: entity work.fofb_amp_entity_8b25d4b0b6
    port map (
      ce_1 => ce_1_sg_x92,
      ce_1120 => ce_1120_sg_x32,
      ce_2240 => ce_2240_sg_x28,
      ce_logic_1 => ce_logic_1_sg_x20,
      ch_in0 => register3_q_net_x15,
      ch_in1 => register3_q_net_x16,
      clk_1 => clk_1_sg_x92,
      clk_1120 => clk_1120_sg_x32,
      clk_2240 => clk_2240_sg_x28,
      i_in0 => register4_q_net_x14,
      i_in1 => register4_q_net_x15,
      q_in0 => register5_q_net_x11,
      q_in1 => register5_q_net_x15,
      amp_out0 => down_sample2_q_net_x20,
      amp_out1 => down_sample1_q_net_x20,
      amp_out2 => down_sample2_q_net_x21,
      amp_out3 => down_sample1_q_net_x21,
      fofb_amp0 => fofb_amp_ch1_o_net,
      fofb_amp0_x0 => fofb_amp_ch0_o_net,
      fofb_amp0_x1 => fofb_pha_ch1_o_net,
      fofb_amp0_x2 => fofb_pha_ch0_o_net,
      fofb_amp0_x3 => fofb_decim_ch1_i_o_net,
      fofb_amp0_x4 => fofb_decim_ch0_i_o_net,
      fofb_amp0_x5 => fofb_decim_ch1_q_o_net,
      fofb_amp0_x6 => fofb_decim_ch0_q_o_net,
      fofb_amp0_x7 => cic_fofb_q_01_missing_o_net,
      fofb_amp1 => fofb_amp_ch3_o_net,
      fofb_amp1_x0 => fofb_amp_ch2_o_net,
      fofb_amp1_x1 => fofb_pha_ch3_o_net,
      fofb_amp1_x2 => fofb_pha_ch2_o_net,
      fofb_amp1_x3 => fofb_decim_ch3_i_o_net,
      fofb_amp1_x4 => fofb_decim_ch2_i_o_net,
      fofb_amp1_x5 => fofb_decim_ch3_q_o_net,
      fofb_amp1_x6 => fofb_decim_ch2_q_o_net,
      fofb_amp1_x7 => cic_fofb_q_23_missing_o_net
    );

  k_fofb_mult3_697accc8e2: entity work.k_fofb_mult3_entity_697accc8e2
    port map (
      ce_2 => ce_2_sg_x38,
      ce_2240 => ce_2240_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_2240 => clk_2240_sg_x28,
      in1 => assert5_dout_net_x1,
      in2 => kx_i_net,
      vld_in => assert10_dout_net_x1,
      out1 => x_fofb_o_net,
      vld_out => x_fofb_valid_o_net
    );

  k_fofb_mult4_102b49a84e: entity work.k_fofb_mult3_entity_697accc8e2
    port map (
      ce_2 => ce_2_sg_x38,
      ce_2240 => ce_2240_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_2240 => clk_2240_sg_x28,
      in1 => dout_down_x1,
      in2 => ky_i_net,
      vld_in => valid_ds_down_x1,
      out1 => y_fofb_o_net,
      vld_out => y_fofb_valid_o_net
    );

  k_fofb_mult5_ed47def699: entity work.k_fofb_mult3_entity_697accc8e2
    port map (
      ce_2 => ce_2_sg_x38,
      ce_2240 => ce_2240_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_2240 => clk_2240_sg_x28,
      in1 => assert8_dout_net_x1,
      in2 => kx_i_net,
      vld_in => assert9_dout_net_x1,
      out1 => q_fofb_o_net,
      vld_out => q_fofb_valid_o_net
    );

  k_monit_1_mult2_30ad492eba: entity work.k_monit_1_mult_entity_016885a3ac
    port map (
      ce_2 => ce_2_sg_x38,
      ce_224000000 => ce_224000000_sg_x7,
      clk_2 => clk_2_sg_x38,
      clk_224000000 => clk_224000000_sg_x7,
      in1 => reinterpret1_output_port_net_x1,
      in2 => ky_i_net,
      vld_in => ufix_to_bool1_dout_net_x1,
      out1 => y_monit_1_o_net,
      vld_out => y_monit_1_valid_o_net
    );

  k_monit_1_mult6_71da64dfef: entity work.k_monit_1_mult_entity_016885a3ac
    port map (
      ce_2 => ce_2_sg_x38,
      ce_224000000 => ce_224000000_sg_x7,
      clk_2 => clk_2_sg_x38,
      clk_224000000 => clk_224000000_sg_x7,
      in1 => reinterpret2_output_port_net_x1,
      in2 => kx_i_net,
      vld_in => ufix_to_bool2_dout_net_x1,
      out1 => q_monit_1_o_net,
      vld_out => q_monit_1_valid_o_net
    );

  k_monit_1_mult_016885a3ac: entity work.k_monit_1_mult_entity_016885a3ac
    port map (
      ce_2 => ce_2_sg_x38,
      ce_224000000 => ce_224000000_sg_x7,
      clk_2 => clk_2_sg_x38,
      clk_224000000 => clk_224000000_sg_x7,
      in1 => reinterpret3_output_port_net_x1,
      in2 => kx_i_net,
      vld_in => ufix_to_bool_dout_net_x1,
      out1 => x_monit_1_o_net,
      vld_out => x_monit_1_valid_o_net
    );

  k_monit_mult3_8a778fb5f4: entity work.k_monit_mult3_entity_8a778fb5f4
    port map (
      ce_2 => ce_2_sg_x38,
      ce_22400000 => ce_22400000_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_22400000 => clk_22400000_sg_x28,
      in1 => assert11_dout_net_x2,
      in2 => kx_i_net,
      vld_in => assert12_dout_net_x2,
      out1 => x_monit_o_net,
      vld_out => x_monit_valid_o_net
    );

  k_monit_mult4_1b07b5102a: entity work.k_monit_mult3_entity_8a778fb5f4
    port map (
      ce_2 => ce_2_sg_x38,
      ce_22400000 => ce_22400000_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_22400000 => clk_22400000_sg_x28,
      in1 => dout_down_x2,
      in2 => ky_i_net,
      vld_in => valid_ds_down_x2,
      out1 => y_monit_o_net,
      vld_out => y_monit_valid_o_net
    );

  k_monit_mult5_a064f6aaae: entity work.k_monit_mult3_entity_8a778fb5f4
    port map (
      ce_2 => ce_2_sg_x38,
      ce_22400000 => ce_22400000_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_22400000 => clk_22400000_sg_x28,
      in1 => assert4_dout_net_x1,
      in2 => kx_i_net,
      vld_in => assert9_dout_net_x2,
      out1 => q_monit_o_net,
      vld_out => q_monit_valid_o_net
    );

  k_tbt_mult1_cebfa469e3: entity work.k_tbt_mult_entity_b8fafff255
    port map (
      ce_2 => ce_2_sg_x38,
      ce_70 => ce_70_sg_x27,
      clk_2 => clk_2_sg_x38,
      clk_70 => clk_70_sg_x27,
      in1 => dout_down_x3,
      in2 => ky_i_net,
      vld_in => valid_ds_down_x3,
      out1 => y_tbt_o_net,
      vld_out => y_tbt_valid_o_net
    );

  k_tbt_mult2_2b721a52a5: entity work.k_tbt_mult_entity_b8fafff255
    port map (
      ce_2 => ce_2_sg_x38,
      ce_70 => ce_70_sg_x27,
      clk_2 => clk_2_sg_x38,
      clk_70 => clk_70_sg_x27,
      in1 => assert8_dout_net_x2,
      in2 => kx_i_net,
      vld_in => assert9_dout_net_x3,
      out1 => q_tbt_o_net,
      vld_out => q_tbt_valid_o_net
    );

  k_tbt_mult_b8fafff255: entity work.k_tbt_mult_entity_b8fafff255
    port map (
      ce_2 => ce_2_sg_x38,
      ce_70 => ce_70_sg_x27,
      clk_2 => clk_2_sg_x38,
      clk_70 => clk_70_sg_x27,
      in1 => assert5_dout_net_x3,
      in2 => kx_i_net,
      vld_in => assert10_dout_net_x3,
      out1 => x_tbt_o_net,
      vld_out => x_tbt_valid_o_net
    );

  ksum_fofb_mult4_ac3ed97096: entity work.ksum_fofb_mult4_entity_ac3ed97096
    port map (
      ce_2 => ce_2_sg_x38,
      ce_2240 => ce_2240_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_2240 => clk_2240_sg_x28,
      in1 => assert11_dout_net_x1,
      in2 => ksum_i_net,
      vld_in => assert12_dout_net_x1,
      out1 => sum_fofb_o_net,
      vld_out => sum_fofb_valid_o_net
    );

  ksum_monit_1_mult1_c66dc07078: entity work.ksum_monit_1_mult1_entity_c66dc07078
    port map (
      ce_2 => ce_2_sg_x38,
      ce_224000000 => ce_224000000_sg_x7,
      clk_2 => clk_2_sg_x38,
      clk_224000000 => clk_224000000_sg_x7,
      in1 => reinterpret4_output_port_net_x1,
      in2 => ksum_i_net,
      vld_in => ufix_to_bool3_dout_net_x1,
      out1 => sum_monit_1_o_net,
      vld_out => sum_monit_1_valid_o_net
    );

  ksum_monit_mult2_31877b6d2b: entity work.ksum_monit_mult2_entity_31877b6d2b
    port map (
      ce_2 => ce_2_sg_x38,
      ce_22400000 => ce_22400000_sg_x28,
      clk_2 => clk_2_sg_x38,
      clk_22400000 => clk_22400000_sg_x28,
      in1 => assert5_dout_net_x2,
      in2 => ksum_i_net,
      vld_in => assert10_dout_net_x2,
      out1 => sum_monit_o_net,
      vld_out => sum_monit_valid_o_net
    );

  ksum_tbt_mult3_e0be30d675: entity work.ksum_tbt_mult3_entity_e0be30d675
    port map (
      ce_2 => ce_2_sg_x38,
      ce_70 => ce_70_sg_x27,
      clk_2 => clk_2_sg_x38,
      clk_70 => clk_70_sg_x27,
      in1 => assert11_dout_net_x3,
      in2 => ksum_i_net,
      vld_in => assert12_dout_net_x3,
      out1 => sum_tbt_o_net,
      vld_out => sum_tbt_valid_o_net
    );

  mixer_a1cd828545: entity work.mixer_entity_a1cd828545
    port map (
      ce_1 => ce_1_sg_x92,
      ce_2 => ce_2_sg_x38,
      ch_in0 => register1_q_net_x6,
      ch_in1 => register1_q_net_x7,
      clk_1 => clk_1_sg_x92,
      clk_2 => clk_2_sg_x38,
      dds_cosine_0 => register_q_net_x12,
      dds_cosine_1 => register_q_net_x14,
      dds_msine_0 => register_q_net_x13,
      dds_msine_1 => register_q_net_x15,
      dds_valid_0 => constant15_op_net_x1,
      dds_valid_1 => constant3_op_net_x1,
      din0 => register_q_net_x31,
      din1 => register_q_net_x32,
      ch_out0 => register3_q_net_x15,
      ch_out1 => register3_q_net_x16,
      i_out0 => register4_q_net_x14,
      i_out1 => register4_q_net_x15,
      q_out0 => register5_q_net_x11,
      q_out1 => register5_q_net_x15,
      tddm_mixer => mix_ch1_i_o_net,
      tddm_mixer_x0 => mix_ch0_i_o_net,
      tddm_mixer_x1 => mix_ch1_q_o_net,
      tddm_mixer_x2 => mix_ch0_q_o_net,
      tddm_mixer_x3 => mix_ch3_i_o_net,
      tddm_mixer_x4 => mix_ch2_i_o_net,
      tddm_mixer_x5 => mix_ch3_q_o_net,
      tddm_mixer_x6 => mix_ch2_q_o_net
    );

  monit_amp_44da74e268: entity work.monit_amp_entity_44da74e268
    port map (
      ce_1 => ce_1_sg_x92,
      ce_1400000 => ce_1400000_sg_x3,
      ce_22400000 => ce_22400000_sg_x28,
      ce_2800000 => ce_2800000_sg_x4,
      ce_560 => ce_560_sg_x3,
      ce_5600000 => ce_5600000_sg_x12,
      ce_logic_1400000 => ce_logic_1400000_sg_x2,
      ce_logic_2800000 => ce_logic_2800000_sg_x2,
      ce_logic_560 => ce_logic_560_sg_x3,
      ch_in => ch_out_x2,
      clk_1 => clk_1_sg_x92,
      clk_1400000 => clk_1400000_sg_x3,
      clk_22400000 => clk_22400000_sg_x28,
      clk_2800000 => clk_2800000_sg_x4,
      clk_560 => clk_560_sg_x3,
      clk_5600000 => clk_5600000_sg_x12,
      din => dout_x2,
      amp_out0 => down_sample2_q_net_x5,
      amp_out1 => down_sample1_q_net_x5,
      amp_out2 => down_sample3_q_net_x5,
      amp_out3 => down_sample4_q_net_x5,
      monit_amp_c => monit_amp_ch1_o_net,
      monit_amp_c_x0 => monit_amp_ch0_o_net,
      monit_amp_c_x1 => monit_amp_ch2_o_net,
      monit_amp_c_x2 => monit_amp_ch3_o_net,
      monit_amp_c_x3 => monit_cfir_incorrect_o_net,
      monit_amp_c_x4 => monit_cic_unexpected_o_net,
      monit_amp_c_x5 => monit_pfir_incorrect_o_net
    );

  monit_pos_1_522c8cf08d: entity work.monit_pos_1_entity_522c8cf08d
    port map (
      ce_1 => ce_1_sg_x92,
      ce_224000000 => ce_224000000_sg_x7,
      ce_5600000 => ce_5600000_sg_x12,
      ce_56000000 => ce_56000000_sg_x5,
      ce_logic_5600000 => ce_logic_5600000_sg_x2,
      ch_in => down_sample_q_net_x3,
      clk_1 => clk_1_sg_x92,
      clk_224000000 => clk_224000000_sg_x7,
      clk_5600000 => clk_5600000_sg_x12,
      clk_56000000 => clk_56000000_sg_x5,
      din => reinterpret5_output_port_net_x1,
      monit_1_pos_q => reinterpret2_output_port_net_x1,
      monit_1_pos_x => reinterpret3_output_port_net_x1,
      monit_1_pos_y => reinterpret1_output_port_net_x1,
      monit_1_sum => reinterpret4_output_port_net_x1,
      monit_1_vld_q => ufix_to_bool2_dout_net_x1,
      monit_1_vld_sum => ufix_to_bool3_dout_net_x1,
      monit_1_vld_x => ufix_to_bool_dout_net_x1,
      monit_1_vld_y => ufix_to_bool1_dout_net_x1,
      monit_pos_1_c_x0 => monit_pos_1_incorrect_o_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_2_sg_x38,
      clk => clk_2_sg_x38,
      d => adc_ch1_i_net,
      en => "1",
      rst => "0",
      q => adc_ch1_dbg_data_o_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_2_sg_x38,
      clk => clk_2_sg_x38,
      d => adc_ch2_i_net,
      en => "1",
      rst => "0",
      q => adc_ch2_dbg_data_o_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_2_sg_x38,
      clk => clk_2_sg_x38,
      d => adc_ch3_i_net,
      en => "1",
      rst => "0",
      q => adc_ch3_dbg_data_o_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_2_sg_x38,
      clk => clk_2_sg_x38,
      d => adc_ch0_i_net,
      en => "1",
      rst => "0",
      q => adc_ch0_dbg_data_o_net
    );

  reinterpret1: entity work.reinterpret_c3c0e847be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => assert11_dout_net_x2,
      output_port => reinterpret1_output_port_net
    );

  reinterpret2: entity work.reinterpret_c3c0e847be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => dout_down_x2,
      output_port => reinterpret2_output_port_net
    );

  reinterpret3: entity work.reinterpret_c3c0e847be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => assert4_dout_net_x1,
      output_port => reinterpret3_output_port_net
    );

  reinterpret4: entity work.reinterpret_c3c0e847be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => assert5_dout_net_x2,
      output_port => reinterpret4_output_port_net
    );

  tbt_amp_cbd277bb0c: entity work.tbt_amp_entity_cbd277bb0c
    port map (
      ce_1 => ce_1_sg_x92,
      ce_35 => ce_35_sg_x22,
      ce_70 => ce_70_sg_x27,
      ce_logic_1 => ce_logic_1_sg_x20,
      ch_in0 => register3_q_net_x15,
      ch_in1 => register3_q_net_x16,
      clk_1 => clk_1_sg_x92,
      clk_35 => clk_35_sg_x22,
      clk_70 => clk_70_sg_x27,
      i_in0 => register4_q_net_x14,
      i_in1 => register4_q_net_x15,
      q_in0 => register5_q_net_x11,
      q_in1 => register5_q_net_x15,
      amp_out0 => down_sample2_q_net_x34,
      amp_out1 => down_sample1_q_net_x34,
      amp_out2 => down_sample2_q_net_x35,
      amp_out3 => down_sample1_q_net_x35,
      tbt_amp0 => tbt_amp_ch1_o_net,
      tbt_amp0_x0 => tbt_amp_ch0_o_net,
      tbt_amp0_x1 => tbt_pha_ch1_o_net,
      tbt_amp0_x2 => tbt_pha_ch0_o_net,
      tbt_amp0_x3 => tbt_decim_ch01_incorrect_o_net,
      tbt_amp0_x4 => tbt_decim_ch1_i_o_net,
      tbt_amp0_x5 => tbt_decim_ch0_i_o_net,
      tbt_amp0_x6 => tbt_decim_ch1_q_o_net,
      tbt_amp0_x7 => tbt_decim_ch0_q_o_net,
      tbt_amp1 => tbt_amp_ch3_o_net,
      tbt_amp1_x0 => tbt_amp_ch2_o_net,
      tbt_amp1_x1 => tbt_pha_ch3_o_net,
      tbt_amp1_x2 => tbt_pha_ch2_o_net,
      tbt_amp1_x3 => tbt_decim_ch23_incorrect_o_net,
      tbt_amp1_x4 => tbt_decim_ch3_i_o_net,
      tbt_amp1_x5 => tbt_decim_ch2_i_o_net,
      tbt_amp1_x6 => tbt_decim_ch3_q_o_net,
      tbt_amp1_x7 => tbt_decim_ch2_q_o_net
    );

  tdm_mix_54ce67e6e8: entity work.tdm_mix_entity_54ce67e6e8
    port map (
      ce_1 => ce_1_sg_x92,
      ce_2 => ce_2_sg_x38,
      ce_logic_1 => ce_logic_1_sg_x20,
      clk_1 => clk_1_sg_x92,
      clk_2 => clk_2_sg_x38,
      din_ch0 => bpf_ch0_o_net,
      din_ch1 => bpf_ch1_o_net,
      din_ch2 => bpf_ch2_o_net,
      din_ch3 => bpf_ch3_o_net,
      ch_out0 => register1_q_net_x6,
      ch_out1 => register1_q_net_x7,
      dout0 => register_q_net_x31,
      dout1 => register_q_net_x32
    );

  tdm_monit_1_746ecf54b0: entity work.tdm_monit_1_entity_746ecf54b0
    port map (
      ce_1 => ce_1_sg_x92,
      ce_22400000 => ce_22400000_sg_x28,
      ce_2500 => ce_2500_sg_x3,
      ce_5600000 => ce_5600000_sg_x12,
      ce_logic_5600000 => ce_logic_5600000_sg_x2,
      clk_1 => clk_1_sg_x92,
      clk_22400000 => clk_22400000_sg_x28,
      clk_2500 => clk_2500_sg_x3,
      clk_5600000 => clk_5600000_sg_x12,
      din_ch0 => concat_y_net_x0,
      din_ch1 => concat1_y_net_x0,
      din_ch2 => concat2_y_net_x0,
      din_ch3 => concat3_y_net_x0,
      rst => constant11_op_net_x0,
      ch_out => down_sample_q_net_x3,
      dout => down_sample_q_net_x4
    );

  tdm_monit_6e38292ecb: entity work.tdm_monit_entity_6e38292ecb
    port map (
      ce_1 => ce_1_sg_x92,
      ce_2240 => ce_2240_sg_x28,
      ce_560 => ce_560_sg_x3,
      ce_logic_560 => ce_logic_560_sg_x3,
      clk_1 => clk_1_sg_x92,
      clk_2240 => clk_2240_sg_x28,
      clk_560 => clk_560_sg_x3,
      din_ch0 => down_sample2_q_net_x20,
      din_ch1 => down_sample1_q_net_x20,
      din_ch2 => down_sample2_q_net_x21,
      din_ch3 => down_sample1_q_net_x21,
      rst => constant10_op_net_x0,
      ch_out => ch_out_x2,
      dout => dout_x2
    );

end structural;
