`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VMrHUJ7jR2a4on8XaeYhAjIaz4rRbGfwW8VHamgJPReOlpXR5SnSuFHyXpuBXjJtExIdI4sljp69
+hXbGMBP6w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V60B8mHqwCWcAQivsECFj998ByvDjB+8JeAAOvVLZEni4XD/2U9vfLmYo3cbFA7NMwmRaGCTY/HS
60s+TT01wMgHgujfEF49/mRJ1glpwP7EhB84g1K7xdtpOxYzMggfDKm9YDHGdz17ha5r9njnY1zy
JipFw5giX28n8uHL9G8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GKYRZjR/TFpnasPz3c3jVHgchRKQZzQmbeBlvkY7oOgwxypd/dr4VwpVMi0c/+LrTgTuOuMQWz2+
vRSLHWdQymehN5n+43A7V/DOnpsZhWNbBZjAAuoAfwm2rYmgABKSNALo8Z848RWnPvSJMnRNGZpC
9BkLlvkk/FGaUYmfKejiN/kDk7F+OC0xZKM06r67ElLn3O2SM3TuNkYTyDXfz95kCBzmkR6aRsXS
coxZYmkVs3Bzvl7yGV7eK4o+z/3pK18wgBXBXKPtKxy0OidDULBiGLl1ZKQMbtBMZsj4eKSkFDOv
DgdJpMEyup8XzH4YzfI4QinCaVxQwuGZ6+xZlQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pXvJEU59cRATVhmRJ1vsVWJPmFqdKz9UXT5pm7AP0hDS5zf02+kgpTD6arJVkG/T6Lh+I5bkhqT2
BXrjBzlv9yK8zwQamfQphBZUgyovPxbNO/0apAj/dwXgXToNeC8wjGMKOoPVkEAFgLXC9pbMEfXH
q7zz+PYXcMJbejWqEF8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r5I5r1xSDgVITJSqT9zg4YQgFLAtqfFW7eaJ/VcLwoK4wHV3PLEhK/YA8kF7MbXjDSnIB1jq/Lbq
d6Uuvb7kijHkFrESXiLB+MGWUasIWXJUZK9t7gT8tA9FiSeXPGQ83fgMtOifSov62C3dAsdSYWXH
CA2noMSeo1xFTmVQKw81KxLnv6RExz75rRcPSDjnLnjq0wC4qY6irtnNTR2Ksvj6OlRXYQSC0Lnn
tUsCjZyHrR7WdazpAChMTAv7/FNpfqV7Vn+ftdwOXXzoTOyvsuJ3L0sdwjtiFmDB7P1LM/g5nIHl
nUJ408y1B08faieNRdh1D4XkCbRg017ZqjwE2w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13392)
`protect data_block
KtAu6lOpfhhiJMKUeQgWfQaqAFeGT6VM8dflx+KL4IWP22gxzGk7dVp3rYdTkOJTcBl3oC1L91cx
/1Cnv0TE5rO1BXSRtTIlnC62+xpU4iNdOsPkWXJt4ImOpV6V3uck6luHN0ec4jQwmhLTx07XSPmD
VO9Uj129zbM2Sf57PVGBpe7nbK79iv9e8bWeo0ekO1kEqLRejlsK9sjxoxM8dcXpXACbpn5xJ6c0
p4i741eSxyKHu0ejKMdlMoTDjvmWAaW4oUQMPKwaRBDj6TdjPcBIMqqdbjh0HoPRYO9MzRXdNoj/
IYQsrXWYPACKFPSWeFyk+SBkA3ZU76pLIhasSm/sttOri9EBG16/6E8Z54aRpnjjYQsutIIM8R2j
Hdlzz3lCRMIXZdEaNnODfv5Bs6PqEBLhpWFiMsLM+i+jlRoyuHJ6xjY76w/GiXXNenaqyYIR+APo
RCcXaYdqFvLDm1p0wJvANDawiBdRVxwj1xLbzveQOt3Ln/s+dgCbbr2ktQx/XYCTkzNrf1DojRQs
DpZ+FCTYDM1W2+XVHrgMCccLMRcH3QgUvZLdMv1UtqmPuzbyaDmLJaGgrNFD2wLdhWv1pPsPiGTV
A+PICqpCnuLCD6dvuuDYfiE41iifFzSWen1OZ92DZLCzdnq+NghuPPdg5jAW/ajyq42scJ783D0a
2K3s93M2B+flxrfpvB9RVAYqDXg7ekpuBg+rPqDicLSOULbmHEr5nEKWoJalwLEvH5fXuLWNfgyb
/Z2xtHnRJTerjPQHd4OdB647tIYVcn+FCg91U5NC3Il+CEKSWYln0HQMvu1gK0vWNaGldZvsJXS1
ER2WR+woHT5+uocyWj/wRPjvHSFPyuE2VzRV1GdPYshxcMkFi5l+kWXpjadQuZVTViigRb8Z29GA
tj1kB67Y2SfrjRLOuOZVTW6PhByEPMnfp4iuupAL6OM9+IYOLkqmytw3hn3TxZz6w1rSojvRQ6V2
JTiFdIevPwCi4kSMf9D0e9+vesa+g0zACQur0GfGrnNtkgn/N65WqV3HQT04C/lc0T8KXRXHotv2
KR0E2S/U8c+YmqfamQ5kFNBnQnwv4mPOU6ETVMiS2YWoDLjCkwUbRTK0nvdVDMItW5PWrGAwqPLk
x8lrqCk1HWsRqqkJr6aNPxPOHvMTOqXgvvaXRnKFWnyc06YpG4Wi7Wz1DkDCFBpCuzSI4K3WJA91
fmSuK10HtfLQzETj6QBCDJM8UHaSi1KBI+lZEX3O8tDiNonS/gJkf0KuLt4Gg6+ZO8/WWsJtd+Yo
Y/MCM6gG10i5qOohsDv16MoM6c91u5uwvXsavqfjuCy4JFa+RdANwf1NmmiYf8yxBi4foKqWBvlu
XQuPggLbGzAo45Z45T/Y4oBUZSpRa1FwunUxJEnY6RjLhxkvUbOf6FFgPa3TVqw752urFFAb+RsH
S8EgIeawlQH2rmTOhEJBfJRb16zQ/3xaLiS/6kLsE5JBqtgrb3mKVqh9PCyWOmseHT1AxBr0+aP0
GBG/PyBaqfgIk+9fIkW2W1BTAaz04eDtv3cF5m45gg+wzKTckS8BNk/+tTEhv+hQgQxbdODlqofx
vrZto4baZaHD+M7V+H59TENSaGnzd0fXJ13MxG29qoXrCaJ5HlPT9n09WE/9WC/sOC60PHos3B6G
v8Egt47JBvrmDcgljBvYHnxOFVmLXwx3V5tFShRUmq0uGpbibXbTMkxyJURlkJCc+sXHp6bh/hNh
XDJCesEXQnuWBUk3lhyc2LdgXhBQDjsl5ezP6s0UqE5VXe0MZS8Xu6Y93WP4ApK4fMUcKBqjfxU7
gx+F0zEXX/tUOTchTPLZXCC/R73+ehq6ZSKjIo/PsVkII7G+G4zC6tLCa8cMFSua1Egi7VaRrv7h
eOX2SgKkjboJK3H6DoqdH5sUsAgsckWtj6EmADCfWgJPJkziQYD2X7hPEpxU69AHBw21bYYCdkE0
L2sbor15Cet6k8wZmU5Qd9AdDa0rzGP2vQwCQZfy8xfOnkCExm4keLdGvOxedFkX6oCou/OZtLC5
seQDxm2qdyV9tmKrUlZUv5c2EE8PiTxhVnCXeU3EA0Fsy7YFXR9KTSqZJVOhSvbu1834E7v65yis
+YgdquOItIB/dujyMKyWMHsxkwtGm3/nNpW7SoYyqf59qTefO8gcOFwjujLMGaX8xLx0bgkG7OKy
qlCAZl02XYrHsXSe7OpYO5NAdu5nKR17+QDG6uqMNdiItPXzZxH5M6fVZA9gdmcwKsI9iE3+a8Vi
/fNq5/wTd0ReYWEsueU0YKFbvNNgLf/dqPdylVuU8PKhJrHalElU62RDyLfr724GuhBdGDBlGjoN
1UdE3fe+UzcUQm+fRi0JDByqI/H/yGZgWAmE7MY4thSx8HkJf6nMRjr8u4SEjwix2IJ7Z5xJpQGF
qximcuXUIk6cX1FjBq5Sd+Ozk2JmWvxLfA5uRjeJwRd109thPcsQ3gEZG6Bm1wfr7W/ZpKD+1BKL
xMSG3jj9cb2pxmn7D3Rah3q1TV98H7T8sKN9h2j2ZaytJNU+ZdHG80ZKkFVMDN3m1jBWo93SkqMn
XnPSsVVBAkvy1NteShwmVUKh1HI03rG8ORyOs4zEcygSe9NWnZs6ytiFaxChj7sjzYdJy8qaVMtf
enFAkp9VtCM/YL5crMVf5858JuM4l7tTXw9DuxuddYI6uuz4Uy5bTymZEASwa1/+QnSGXkFyfjQe
E4SqVO2VcPiZ2TA6CHFTM4gMVoC2w954suZ4YRP2Q4h1X77cZlIo9q7ZESFPneNyg9TteU4+cl0F
+ZuXnhUGRTtWZQKD3mkBQjRBytkgXcZD/AEm+E5kFRQ4gqyK2UjBm3x4ulu4V2+kqZQfUVVXVCPB
pw5EwMMqB6xfbu0N3YZM6Pj8Y9l8zORPdp5AWioiHByEdEnm6K4tGx0Wzd7vCfUoTmZdXlCa7vnA
dCOo4VSrpw3tijA7Otl7JtVe1HcIYzeCGzsYhzWfGgKeO6J3xxJSWqSXJss5c72gctvTkDGJ7L8m
KyfuFVy1BA1Os9QxrRdLPiuptc1EGnHCQB/Z/3t0JXQ2AAJwWWE7EvPIGoBA7C0XSM+IPCC4Rp8u
F5eQyIjJyp/3Xacg+A0M36sZjQ9Tv0ua768/q1xufC7MUYxlPlr/59mxdSXhCZoxQyAzq0ob7YA6
GfG3HhxQ5V0nlJdmdN3rtyQZF/x2Mb4BABO6pXgrP+fyrzlZtVJI7ULGEWRp4O3Cke3A6h6RtVXk
Kal75VSX4fguegatIjvj1QMwLlyr1s0Ehf87ADEE2CiqordMZWZABgbApTrI5MZcSLpV7ixon0BC
z/zpFPcbPPPPzJ1kBSq9f7+POuEpo2qfpnqe4nKMDiCNpJA1XZc9icX0gcNpaMD7pLAFZmYnOZWI
HUxZ31aWnkwzRExkUbngQKPbXhsBqaBiMufzC/cA6iXyNataSvNI475Bx/RdxiTukZezLR056F7H
bkNQ6IiQyhzJMvOc4Fy1Ge2zDtZOffcD4FKL4b9pEPJp2MLZB4c7dwkoK2zFj0/6O6x+uaeCj/51
UnlP9k9K1O/Ek/y4Q3D3xzvuFxLwX1E0hbfe4dDgsMQPfD6LPY5A/0ZLGxTzYC3gxuiP2tnM8BHm
xqFmWmIGL8Nkj5mLtsOwURE8fdksfCw6HGRj4nysOmK/D9tA2LaXMaKu0tvab0hUbxnW/DUm10UI
RR4PyIHO+66KjYapXAalXWBw6bGR9uiOUuzfP0jzD/j7DfUEznFuGpYAkfxtHZbSKERWzVUlQEhi
uwyticDxBg5o7mkEQnHuREykNRAbz9OlqUdtpzk/nbgDtcCNuF0v9FHk/EDe3wzrX/Tj98fcRsRf
aAsyPb6nIG89ioTWL6ZNmxF/Ft0ma6+liPBqGaZ7pG59gyvzMIujhLP27qlbWvqtxwd5IW69yfJc
Rpd/bSGQKYpRJrpHN3hGIdsyYCyuyB8WIGeaElRlgZwBE7eZI5j3GlnYjGiefE4eWJ+CuAkQnvyO
yEQfbERrLSpEEFS9oygelpLIWtIUfa2+bypsEilA4ccH3ALJhnbOFguPlGLpJs7NlexiJa9xttgA
tWUq22F0Vl5Cj1kZvtxGZMIfQCwSiYMS+daS9PHhtkqrylJtsbOTxYEhC6dO+v79rr7LH5UMLuhO
Z3KrJ+IVdwlOA7sexF/1duCreNLBbnYrp+VPnJCK1LpPfgtSlWk+/4wHEwnLmCysbO6TqeMOX6z8
RFYv7o+GN9XC756ctoI4aFVXWhltwJVUrcr5qqK7FZ6xLGhjdVo2VOEQWz/bc9qM1u2teBRzOQIk
ksCQcPrge/Zni8HuaEqtP/8mx44KGlxNUhFJW/eNrich/lIBLOt7JqDRc89+TK60q/W46arZ+BEL
IbOukqGcixAht4NtdA8KBJLac72folUZFyq6uMY5SIpakCk5puD+jLYwzGfciJzGzrLInKiB5lzh
V40TUVUfZMccYoeOXHdk3+T/vHthMO9nZ2UIWApEUdusSYRH27Dqvk0eZXxedBXtHBJPhxxIiZ8p
EbpwXKmGXVGMQIbY75L3EbP9Y0LNK0so9CYZqivll+pUKOpyLOsqDGFdG9ayqwy7w9J6la/W8h/h
fCZmzHsUFLCrHXyF5p9r8AL9GGdc7ReIZ9sNdAlfOxI/ZEx/hbnv7HFDrBz3Xx117NL0DvNzMBcf
Fiazfjgk3tthUkGiFgIyjy25PaA/k52kLIq4MAyIFu7O2dZuiyD77jjAkZG0hK/om08L2Nq9+wpX
wY6m0TnwDLggEqT+ojgeSh6gI72AIZvnRbDRMsR/wlNRQYksbX5yq7cp32CqsYWT+/Rg/jue1Bnc
7wtlBBec9KDMQvgYre0GJ/pZc0wRG0yeOjaUJEgd3Qw9S6jNcGglR73A7TWQ7HCspRJkQYneEdVO
xTls5U3jmqoB/fAJvouUmUEyskQRXzQyPGISIE2ZJLW1HXA9oFQvCcXCJGEuXdixoHU4QJssRgSd
k0OFyC29yVWF8s2LPpjfSi0s2JfrG6tLjN9LkNINfZXe072f3sXdH+XfjwK6erUscc2YxkGiYTWJ
V5E6e22ApEPsEhG7kxspUQi/OB2JDo6Gns+30iUR2y33HJ4ZWy6ttOxrEIlkgKFS05hQn9ooirQL
EbuOeFNbPsGUQ53+Gyz7GZuO3PiWpOEhXvk9U7HfMW0XWV3NEAhnN67vbH7A51I/sgnrkk5W8iL1
PV2vcb6H2TUa3/cFfcnaJSIB3NwP8wvFt5Lu5YUtf59D6mRp/JAutb8FApD+Bz69T22LkrISdxIz
Tk1gern+mDrUuOGu/guIHNnYnR3cY8meDhU1Tw4KgjND8k7bO3XvhUQ4DL8/FERDc3Hu8ZkllG4X
xe+qzUY6Jr4iWjIurCfQQ1yFehXf8AFvO970wYg/W9brH2/tiazw6eMMEH/vGl6pbus4Ydzq+RDa
zRLXrEKb/l0QXkZaK1qr51T+9qoFS1gpQQbwvV3MFfm6oviHkESYHQmr7vBuJMWJgGUYaQYANeuZ
aPFiz8h5lu4j5dDOAGPymmFKy/rjnhRrj1h5dfOfCUjQHkuokoRpfq2hhk8meY1jjT6Mq9KqAhY6
DdGQg+VT7RNE68ZL8/UkxP5QJbpiDVXcMAsEcSdW8g1JLHOazsbJczMEWWrFJFNVG0/QOri3ykni
vNCytio4klf7TBY+JeGNPm8bRifJt5voKJZtACxE8H1cR6+Xi+vvX32+BJ1CjcbUQZlxlBWiopan
2LIXFllhqwR2R4ePyMoCsgsQNqdKPT5rhk4Qu6ZE42DWGKJYijDLKwy6jt2GvX5FvdPC6Zot7QmX
YpaiJxxoVM/KkpBg0ezNJtEyGH0EOOyamVVHtbgyF5+4Fu2rxk+jcwhHxwHneBocmuXt1v/jw/XJ
a/mO+goEY+iV6g7B8wvkF3Gp174s1cm0sIgla4WU8TN1Rhx1K89egoY+NLH88Kr1dLRAaFRI/Ra3
+r/va9E780Z0B6UPXl/wc36fgSfyuwh+0qehPOlsmhyq5CYpVyhfhrTcdfIFwgJh7pQuJpx+wa/C
ZShtqX4+1WA6YtusYrAHStAC8f/COdQvkraoeEaETqrq+k4WQDYNfWFNXxt8N+1/lvi0Q1iOjHSM
Jr+omK7G/y5pgZjmyZQ3Xqv3HhwAX+tJtOBAtywGEwUrzHAKRcD+IGzmwQNE6+Edu8AhclD1jiho
I1TkNUNcr7I8tbN3AgXy9uMN+Xl2576TN51ppNqX5WQBhI6NbdaXvfZojCd9C+n8ZAXaJMXd5Pgk
OHBtILdUfUrXjaIj6UMkdTP1MmRfX2D/IgLUVDoAfa2JURAF+PNoCbNR0/uG2zeuYccRSw9Xxi0T
pm8VimXiGd/w14mqIYtbE9nw52Pe+uuMDavHlP7hMk6ZQasLjI486s8PkkPDvqbvPRi13oWjrA8M
YDoilq7EyDh+krZy49kdeDNRHDOe1YPQFArryMmBEinJsnhvxIc/HKyzbKbz9LYR908id3Aezxmt
c9TXQTAEx3Ju6hvkE2q648++10Yhzsy/9mX8jLrqsVLnKd9M7l23HxkOwgEHAWC6ebjf1pF1ar9d
A60Kq6eX2GkJhcALBa+zzGVAniOrXQYAT9A9w+X6Au4nXovDVo5BMrakexRBEhEzOIyXr3/86qCl
UATvA2qAmEb4RsOHYpUlauWcd2KNBnk+9muZ2Q5X5r9eK2FxTF+1q2RPnP8SCZjgKFsTBQYIDxso
0m9BhxSdWpTK2BOhAPmPYbp02DHkDzyy/0T1TtZCUlwSyGK5P4pNIeWgpaChv67J83mWH/zzxjl2
bRA3BTLW/9UQjo13IMpwxG7fXdjow9M4E0eNXOQJhQapSZbac30rdgJmUsGICbxbsiS0ENB/Sf0w
+/ACabb/y3CUXGHELlWQ9ZjdPISKSPpYhBX4KoiAHo6TECeMADrXPuYQ80mNalKN/OvG1JK0c6Xy
eF02NsfOv4PguZSiZh5zUABkiui/cFvWLD7ZmfTEEQ3Yf4jbBx2jA/j2c2tGo3RjksAjfOIGuOSN
Z9RPfjSpBaya9Nuabbzhax02r7JoGwv7dJBJ/zQb3tx7fPuMAzL/hKoSr+ee9d5ZzAEFpBvMw4Dc
2gqoHCPQ1lJ8Ec/mo+axX3lZrK3WnJ3DRmH/zV217ehNvnAwWag2dzWSeU8WzQ9NUvz/gcw/0Cam
MtKL1yY+TVpxIAIq3RiU6fu4K/Q0k6IHloxasxKwoy+ZiTZTrd6KHQrOZmUc7XC1BeJyzyEnbDUo
ecgDvFCyE/vKUrawJOYM2Wjj9vtidY98UIhgVnewdI0INrcQAm24JmwW+XxaA2VzD63LtPDtGBUn
3NMuSQrLBGvy+XMJU5E4PtA1vSWIct4G/+TPvfxx2Mubv5DQXTIEvVfqSFtQ1exMGhzJbKsTr60V
ETWiyP2quBHeFaevlGfTabbPpu6cmqgAdFCAntS3KHLO2DwW1DvLybrUhBQsPm+b6kDHfFRe0y3J
06Uefsm33g4xCqszeTcuFSz6B75NJsNA7yJZaiVSE8BUFer84bON0fMOc2kaKXw6Khkv+tIHGoCT
t+fzhDK+QposUpIQMZbqOYePQWqB8/uUmqR953z98UjcxwgPeWk2LmTKX5SyMw4WgXRHz8I2TX6k
rhrfZYqy5vuAwsuPxJe/sYxt8PUPf9szN8FUvViRwou/fJErjq/QEVOTEXKRqwE4Z5LPmY/ETzEv
Q+TePW22qr0MnTvD6kk33FAuU9FvvVf9uMwG/izLcM5q1d56WcgMFrEGwS+mqqSFGt7U12AJAASw
Ym/RKudAYH6z9v1c1NOaoRJQlwPm69eJJI7wkAAI6xKOyM+x6/WbddfMS8c8Z3NCDclaimFwvrBT
r5zIs8sBX9M1te7tN7ohb/4Vi/oRilPpbb6BUIC/nyYZOLPn3W6sadcJgTet50R9Ivgum7y2F9nr
qC2aZjqE6MkVTbYA8eJLDsxwsQemYQr3y8beE2xJdPGJurQpirHak0lLatKhYh5j2A6bIrFUA8Sf
baAY2qe5qaEY8Q7fH9LawEW5GjLFGPW/PgfczM0xytXUHmgBRlc9vwKDow1dPtWYKCN2ByrBZQY6
Tb3oAQ565/t8/h1yzwL+HLJp5CXV5gHQyOkXA8DawLgdjaN5Lci5Rr/0BzAOrslDiiuY/j6LoOP+
6LYgR16u8UuSPmpbIGqXpXD6ydxIQ7p51f7v+dg2EMaNwcXBZzvLZIC6sZsgNt9TGkI/2jF22P7X
3XHqTC495EIVuDSowIVkakpnao5uqVJgnhwmziZyZyt/rrBXRa0rZFcOnv/GQlLJQBxZvb9mZbP5
tf9hh5536LpFXnyXsqo6oMDn2biwdRXdKKpc+AZwlhfoCWuzWoGf2c07znwPnyrszVe9quCbirKo
vhd255RWyjLPQG7ZVron0+jNGmqnh5/5384/kpP7u1WIjgCdq7lH5AVjyhnXTBuP7hf4y8e6fGT4
eyhtA6Of/EVP/6pyiikipN41SgrDXJiernEK9l3+P4gR0rLJWQx3QcXEZ3pdo7rIkKpFZMY/6wIT
YPurAqGlKEYR9O54h9NgOmdqUbne/ZzOzfNWAQMZeA+XE/eSLWclD3U6lip75LhN8IVPnfbz+Qb+
aSwAv1ym5mUttYXZ/J9VbKlKCuuJyNE2rlLPJUB4Rhwjwb5tkueu0k2mgw0cAIEy61lNgbntyZ4K
7fAGDpb47IqlqqUqljNBx9m0n9HBNNDpRQTn9a8bTBRALcLyPvXMszwblahQo8HR8gAhKknn+5LV
J2GTKzVFp53GsZ3h63MubwnOq7kurmEjzAJcmfh5gvH/rdGIsn219gZNn/dUNnrmRvRtUmr40eoz
W6diYzOaGHzwUtabGgPrLhQNzQWtmLfIPFBqBHb7trk2FwM38XE2DI6+gEd5wN9GL8mFXXrxoZXU
Wc4+iQjIytprwMm5XcV//J3hUv3GM6zgqPk1e0S9d4L5AVLvsHmTQpGamDGyHBdx93P2X2bi/hCb
HG26sxpiKP7z7koM7gz+2JNXjqjq1lhhlypdztsMpqeK1ymIkzZO9JXJC7W/7h7YHb3Ksdns+GH7
GJXScZDf8SCs/Yb8bUo5581o4fJaItcwdGvZwzqQr1HkvSQwOE/V2bSXXg7vPIv23HZnJibSrMq3
6OBL2OPnaNlFprgIXasrCuesOrJ11E735xQZOLN5YFzy4A0TamHGoTHSpquJ3Pjc1rZ4nJvQU50t
MwRrQYmRPmq7eJ7/zGMgSf2JAc1NTmnJ2NH2qQiY2G/+ofhv17AOk/83tBY6r9wvXz/bZ+2axFui
IsDeWFiB7tRZZ5qsfN7drLVulAFkjnXXLkoedilcAHMQT7pzwTq0KiGStj5cmppNG9rS0VujYXmN
lEH/V/gHtwYhWhCSYBMKzAKgG58riTszrT0hF+C+bmGoLY60ZdFiIIt2qjZX7VUKLSKFGVlmo/e7
pxl0SABnyZ4G2xvVYxvayd/Jnr7dlSi6G1mFJWmcprSoyY6GUhD9MBg5BZ48QaGqvloiUyocE2JH
W8lOE4cf865F0wA9loO4Li7mJEu37cUgGLD1zXqdnrIisNxaigGkJ9PE2ZWMwc6s//8TRLUzM/8T
DDdjcTTG7CZD8wodo3mo6tDjVgXnIPmSArDGUQ0IXLht0M0F5mEogtfGAh7r/lE0lMdjalB4gucG
24u079nF7zZJ3QMflbZ6uRAJTlFeN0BykbP+IcGJ3u6bB4ZNh6E9l6qkZaF1ngNAdeKwtd6aDjgr
Tz6/4fxOj7EUpwu9wfBmZXq8W3aQkozU4r3dXxojXy7RElKYCl9E2Z8JmVJVNqUbp3xBalSw4lGL
WgsBPKzmIFrHR5sp/17fU7A05HYGBqMGzHG6X4DaM7Dw43XBT8M86obHA9oKNEgxqasyXRHkpXRL
P9XBjm0ikBiForWr4wWjr1mMUgjedayKNnswP7RKl7yTMAHuCSp8QWBcv0O5QGxYKMUhmKAAdwKa
6rVQlLA0ycpShEMpHaq4JXeegN5Y0s5/wslzlWd7VWTZNW0UPNYR8jKWHmQ54ul6g3vpotXmQBWE
Fap8RpCzOImagAxXWiu6w51IwhnSh+KRZSfXFmMX7x7x7X8OfnN1lfpSJxusizh9oOg4zbweM+Ek
duOUV1RYYfK8h3ekSyeaIxD3w76zumHRuh93ll97u5irhJ96sQfakmvAaZZbFpoeqGymmof+L3Nh
E0CzucZv0N9ZAzV1dJMz4fpgM+GBsc2Bop+4ukGSyBDF9r7HQd1ykvQf2f7Rhqnb52SbCQKUbYC9
ChG67JsA2Xu8IXrC7NI+ml2UOgsY/+L93o+lJyNojiRh9WZVk5Rq/Zbtof4a3qrmpcIDLGm2fRCD
sXHoh2IQRyIoQtal0hHa7qpje3zVtzhjg4/E9a2Teq31RlsyTaADrvPicr7PAhuczJrrHcSlPL+m
s+0ONCsWcbpNbJJBp8K2i/ynSCqLwcXibJgGTJTN1Ofw3GmLQs9jqLYshfRR05IjYfZRXI63GVNJ
q+0yNYnWfe1JpPhNeJIrcUobcOFRcJwsY/2Y4vteRo+ftk5XyBwT2G5v3xh3mHppyk2w/Tjbr8jB
akTspfi0I8GAMWOQFMGAufEr6Xfq1eQ6XVAEfzjeTD4aklZP3IOqS/XQXu6rb+Qo505z993XUu4O
fjhwhkMgFkspkGXbl3XBQFOKxDz11wmtKRCvj4RE36XFrNK2SEx2y8hp/TzvOKatFsuSeyS+kGx6
q2dFahfNDViA+ClE5lhn2VfkKlkiIrEbvvPOoo1F3DjPnObGqwUkJIfeque0gnNwjXOCN6c5Pu76
pSCtZYzNjb2DQwQhy/Fb4PG8UdDr3xrB03Wsl63+kWschXevY0G9puStYSERw4ayYyFyarcBVY9n
lSuzhMesnDNfHkPTxXcNxt8Z3ryuTrYxETYp0jAsN/ODGLIS5Wr4Bha6QdUeEBHcZRsCdSrFoy01
AhpmWlDsIxVgQKOc+pxkff+rhX+ddDKAnk0Zoq2EuCGgjFFzVaX/LCwuaN6nng1665/yHH9I66pn
RSvM7MdXKNYIXko1COtivHFv7lJvLC18lCTSysSbPI6x8Ld1gFI3wZmKj0PlOgEYUxgDAAy3NdFy
mW2g8oKFJxg8U5ac75GdWE9ook3aUvJX4rb+1vz92HY9wU3SR/3XQGXTyDJeo9iRd9rAS8RY3j7K
zpZ2MNygMUZZhhE1vRjadSAayTRkt9LUgNW2ztdox9yPNL9VCa+2hfya5WvqjXQ2yo2nXZhnNWhI
tHMeSLtDUDfhRxHCgeJfUwlzkBdpaDseRke3BalxinWSTwYjVRirhuQZ+jfU5XZZzxIKz4Wo6OCK
b2MiSMmj1FAHb2R5xnNkKp49jC4X2iv+jSDIOFET8OlmIgXquFsC1AvMJ8403MilqE2owNB7bSAb
1vcPJtt5fc+DMdSTJjj4X2HJzJldgKXz2unLzw0dB/ct4J1pqwc+kBeJESyV//cBKE7aegy1qudR
FohVmw3UtvVMMRc1dcMdaPsA2EoMYgqrjANcyNCiPxYH/1XlYMLmezb65uSBjCYQAqYAawvIOvTe
d0JGkKvOzyJalO5GUjYYQCzTE3vq7j7+gQqEa4yiYx0y7LPzeAn1Z6FEJ0VDb9PY1Q+vTTcQDoTX
vrHPyv3lu+ZhQT1MISgZurCz6eTrIpb1ORRtNnxdIgP8SYFks6FwyzvYZVg7R0GZUpHvPx1x8NF0
VVOCHRSxtwiyjtOG3g2yE7pNq3EMayHqQK2CdtawZT0poUzFtHuHQ3NQZzYDLNTryGKCu10+8Pgb
rzUo6wgy0u4pFiOG3VEeyO9ScdnjPBL+unHGqjRfUlxVIt7hBxexcH9kbXrin2qoq8/eJmJYMqbV
Hc6+uMJohZNssS+N0St1R0Mi6DTZcL/NdEAYSvar8Eq60DcipsouoPtlLq5/yY47E2WxlJpT2uXu
mLOli9Dxcv228mpzKEKK99TDjYwIey/DxMrh9SoQN/s74NbV20Kb2JVe54c/8o2Ml+p5TeCUVQiL
cyzbOCx/bkbYdrTlZhOEj4joVuS2l578uov7UhtiETgHBh4YgxFajCEkgaGx5VvuKkFGYMANuMhk
/nUThEGVwMLI7Bjr8YVE8xqxScKFFF6lRecx2KbELvY2spkFKXKgrkPLkmTZr5rvV1Vp4oKHd+Fu
4t5dEhOQAPOBcmasZNM00Jt79JgAn/uf1ycPmmo2sr9ZpBboFL0hQHk5cYcSC9Q/u2dXUgoeY0Kh
+11b9+4qI5/11HubvsMDGxYLjYGejW5RQfqkkzObfRDuXx1ZRQTYnBFQ6usoiGoJ95xFzxxrg/ir
sO+4X8ytcfn9w7gyM3EucvUUmtvxGeXX+4AHPhmltsvrhC3VyCuY1u56rHUibpMDW7XaAPYshYey
mvD+GLSPyfSkEgRvpYLRA/ZQ3QZuFXpRGE5eBymeoE6zOT8LqELKswR+9/I7RNPXgcPLMsNLkOIX
qB5rLRkzkNzifPfQQYMdhSLlf4D21Ih3SGuLfDMg09BKFvTIWZ3ab+tk1hO7RKtdJVza4vcvL9M5
aFW9W12VmS803EpeRUOeZgBWwJYUWfh0FaJ2vbM6iNVTpv91rOV7eeVF9rKaMSbR7prJjudkhM7L
tQ+aj26ekOjnB676x+Y0p+wBnGX9hEBZ6I+PmY07Q0f8qLE7WgyG42d3OgnDO/4yhTn6Yvk+Fede
EmQl1j+I/LLz/UAuH0QEc/DW623hibsPBLilQDq7wX/hY8S7YU2JehCxtmg1z4vFuqES9fdoI7Kq
Y1TAnXtPuSllLOnHJgWdLPbYEHAh0+QGqN49ScF5xDzC8tuWZWaH50sC4bfKEQPlHLSAFfvdYQ4y
CINNpr5AdBgdtIfTMpsyUMHMjg85PRdWYAiUEpeOi7TgBJSkJRaIO2Q94sk6RviffjzEnQ+RnSLe
Owe+aD5kxhKLH5afl65TnQZfcvH+WKBNhUuQpYN5qdReeTQeq3FiIvl0CE4p5b44ONISt7NictEB
lesqhkuUTpY5ReJ6j4C0Kj7gp7lPWEuLKOA3B2I24tpPOukCrOi0KY9/RpLqWvrTz/x4Moon7+rr
nEtV6FUhd4uFQB05Wzc7w9CAAd6CGdpF00KVGnQxaMRjGvzMEnO2IVPTLz74FFT5tLEUMTauUlmj
jQf4juYyuomuXVRG/y1kv21ZJlDSfhm08LB9Lt/4gl/KcsfTU0zK81hHKc0MkXLvC5zeE7vdKzk/
+xrY1PNmAWYPHa+i/YaEYhRYE0VMOyKpWZHokj1OqVUo4gQa7TV8hDiMqZ0la8csryx1JVhx0u39
lHi+CR8WE8wDde1EK8q7d8p/fvfNSXN16Z0iF+UpayQYtUms03FTZHhrN85296sjdEXE6ZuuQPzY
nvH5yCkGgZBqJoOvP3caqk7i9apKm+0AE4IHCGLdausNBEqduZyMfartesvzzK4rq+7uiqPLLk1b
kT5qGp3+aAHiiWO7oJRMlgdVuFLYbCcDWOllpCoO+XUStIpyC6j2C6PHb4zylWiKQ29T6viOt5oF
D3CjWhcxuUBoNnX7RAJtD255kxVSf4L0viWZE9Mynu/TzHGKPvaezYVx8rCIUNfE7PzzCmUJwxxD
vx4zOLBTeSRgbNPvm4pE8XKCRzJdM6MxrY0mh0b1K3xJnhGGH5dH7Ap5t+iAEeNx9EOnTitWX7y4
r+iHQ+VtqsJOOCOlJ/UZCm2tAVcETx96e47S50XP0RMT8NVVm52sezIFdQ0GpC3gweLVJqWzOY7Y
UeCEwYJE3sHac9DSdHyLxRVhb4H/CUOkKCkW+0KwxrEJAH8QA+B5gmP0BSAIrmlMEbnBV7U+6JTC
gi+9E/S0ZNG5suy4R9vWZgUGMk9eMLKLM8nFTG1/uDxKY/wdsd17pS/+u+IXd1cgp2vi9q8BuAVp
57Uqzbt1jBhAmpnx/0+uRYbN+G9oGUxHhp8jM8UvzQ5kX5vN2R88yzm58ZP1zzjmXYBT9+cfDOqV
+NubtJ/cKHNc61c/9f2zQ1rh6uN6UaPBfhHxJjkBr5XJz/CdxsZi9QydvGZioxGEzCMfARd7wI4F
No/xHuRWtmhG9m9cFIF+0A2PQ3zrVVbdA3fv9n9nt3CPeDiYzFw9qJD84/RJfT0D//YFSEiMzmud
zcsIy8H7hWxTLa9mdh0trPGYzaZX5tdUFz3DdDPEvfwI1mQJfz018dRq1eIaQKKmeMbAxSuCeYdL
lmM5cUJXnEkV1OgxmR2PWgWjuzrDurco/c5BvLJXxEeCVp8MT8mtCKET3g9KHU5z3KZrGoLV3KlR
tzFCehmCjRP7/qmedIa6R61vrt9H90E+Q48vce0Q4XgSmLr2im1ufSqMrLpPP/dejI3sEB7gcwON
uDRT2Ln9X0yFfu0qBAg+rKMDNNgeiInXx4NdZSE5Yqg5sTir0QmS1Rl6lusf/HJFSjx3tQNa9AsI
sJH87wvEbikC9A9QjqLgSv0Bzi2ZQnDfEHM8a0REr9dcGOMlj8C4lnh/vP3jd7fkM6nWT7M/HKzt
dpb2p8VeYEdyocYD1cBy3pv5uvRkViY24TkY5liq/JmAtyAIS4RaPTz0bf19evqcXA6UyDg3ReeK
lhaWn2SeNeqt4otgWrhe85oK7qfjltki1mhkCi5ieKChwJIc7xWc0Cwhjqhszacz1SnFyojlcLqo
4lzuIi2DxoKXuueMZ9bVw4dlfUAbXMw6zfg7g+byAicCnCFuStBznaHSQrQpNSfFW4a40FwBS/I3
+OaUIl9GNGa/frBLjzJWHtkPktwW39e96lbA7+ojFZzaLjLUKvU7M84hYJPem+Tj3w2u1lLk2zVc
5LeQ3QbaWGE0fUKWSaqCLZiyeq8BVQNC4ChmmwhiJU5dFXvF+OGNeecAsSiX5m3+3VSUQUir/+UL
EhGLQc7uhBrtPlANV0oECqHZazsW/RqpOkoddUnd6hxblAGa+QghhJfedzTgTzkflSoUwJkQ0qtQ
QfcQap2AcfUwzzpGWC37cssT3RXms4eWC+BqY+LQnl3rxh7+47RdNGh3c4VdYDKovFuSeKYu5tCI
QOz/6AFOu0lXdIry8DKEZHahrocdkq4YdHSaicurqaW1Zawky87s3Rh/Gz4+NNE/Qii+yBrEk+G4
BLGHj4SX+Ae/lzGqeEplpNmDH0Mz1WBlwSn0IbwqZGBJ3AZhjXSgGK6XSadrloC15slCJdUc8Lmc
3tquRQpDW7w7HMv7BtA93+o46m/HLopQzZCQDtymDrq9DtogHQOIr933uk7hwkA4HxAJq6kpMhFY
r8K46LXLbtB/MfM5TITYP8f7yqt1v4iLwoqY7CcwkVEVoLjqb1D+0tVyhU1L/+mAxgEItELtXhIP
BMjkz4n0PmwqaWLyR16vufaXeBTZ1nvfX4YlaL+nNx3NpmaN5GLiXnIU2o7tAYSDzNtkV5gXgc2J
GlY5lOPw43iH82x2zDOsCgBGiZMXwR7XPA5yk7Mc5CmgXrd7+tXsea6our9orw7KkimoX1bS+8vS
61VEyUwrUDFaG9di6+/z+pYEuGZWnDhF217CEby3QPq/cTZiwBCgCRj8qR5fvuErMWmHPElD/BVB
c9+dogL77HHocVSqE6urXdY4ruVVH8V0I7B+G1KYmxOsySyc8AwFmWcAzhGYCo5fe7iHwq9F8Epw
zeWrEEa7hvDl6eilNRvERnJ0X1d4LEsyq/7Deg7hcL9VfAF+cYG7+tV1aOBJRPngAt7lw/wJeuhE
Rvxii/UyssQ+35HQ4Pnqr+H9pnTbsLP8jCYPeGmXGsYJzD+mxLJyF3DBWQ1XrgxOmF99NNvizLCR
0Y2CxgwGaduANantt60jYQorDZx+4JbCQE6yuy8hIJB7siI1WxTDPpJg1qbV2epgeXMXNyOkzotH
iXqaHpupSqScDQyjtbJYVuys6rvzhbvbvJpiuAYRcxgQsnr1VnG/5kDF6CkX0DOweWd+RsqG9g1u
pNIkVhYvCiB88YkcTPo2l9tkMZRPKyWQ4bgHV+8uVijq1kBz5L5dgc3uRp9gDpC+XZCTdpE79nWx
EEzszvFFj1z6pc4KWzdiLXw0lfEm5AKOhhpwGnTSMf0F13BFWFdWaqx4Jl1gXTny+mO6t2vIYLFP
dPezQUc48hvSGu70A0b7k92tUR8cKkDi3ix5dfaF+kNrH5e/+tZ9ucSbXfID8pu9B6nHY94IWlHG
TuoEESddcDQ8UeMI2doG1f3sUYvRDQhlw4ATWb5jHzGF/2VkOo2FBh6LeDiMN9BQO9nZ4wkeWXEa
BzKjb48bbmXSrfOrOLNY1SGy6bJPRAOXq799/JuI3TWdblnVTpsdLj2xZu+ALQNUHPEtQmCnf7iV
FLIZt7SKlVRl2ut7a2+j+lDi2GXBXgWbvnPFmlcfz4zYysC0Uyq3DMTIKtBEVk51fSUjd2CDlJ+i
s5GrJAEuxFnpwJEgrnH+EMrmKoOP2qwxrtkbaYCijEKgfbnbD11Br/CNF1eLd9DPLepz1mZmSWpy
fQb8e+yUy+PGkL4/j9JOyaKmzB93CFg6tn6EEr0Zfrnd1EZ27nVCcHF1NFEmDpJHeripQEseYI+4
OGkN5cs4ldbMBWInr0JZrYCGf7gQoqkLxsXef+dEJaqX1H9/WTo4Mph8MusECeEcpk+EUQF14aUF
uJrnFdQ4KlyVxz96U62wulMq98JH98/xxifGYGvRgpBQyPJl8U9sT2wEP3kXSustKr2k3ie8asi0
LAI1Pl65vX8KLAlSuAhljxodOdY9/nFoVnc9/irLeuv5sxqFC4/KinqRZoV7PjDl4KwqJ1/t6q/X
YJv93xPSfqq+cjd0JjvY6MrL5PS0E7mugh4Ym4mm4W3g9UZU0FwrswcLyfI19lUA2z8TpA5+ttEP
eFBDuCN0W+Jrv4BNofPQKTMzEFnpExk40LZXtW55jK60lLn75OHCT7pyk+ybbElktUUuVVNtQpwM
+h5CLA6e8zsQxzfjQn5jrXl1do1aHcRzmqaXTPv7zSRpXFITNZHB63ZhOZJJ+AH/5Ta0SijNsEJy
ifwtZgQuEhoKA1nHUlTnFcAqiCxNmxQuIjdtFlwrxnj287ehyR5MY3LPQzKGXwAaAJedHQteMWQv
X0tV3hS/zzFoA6C63cHLC1l2eliJ8zJAFR6/5kEWT3nqzNkTvnXwp+e737psdU9nehVsHg7WAB4e
KDWJQp+eYbY42d+9tDjSvx+nRCVbGMrRIJjbC47R5LaVG0zcASP2ZlebA23CtM3u/Q+LsUH/bp/f
4PQ4rUjY9TamK3cQxmPLumo4FAnzkuK9Uq7sYxTEhoRFP1L+w0ib9M/fcHb7jxTiSQJzzgVo7Sl6
L83NIezjWyGvDEfDaZu01G7bTT0rah4DwqhkPaYynrXOZWXLQfCgEroWQzJtSWE2A/CEq/SY+RXy
qDnO1IYzyReaDt8l3o4meWm5uNpQeoROCCJEGv02qEhWvcN7IvsWgdsy/UVPUE6dgZXc2yLVpC4M
Qy6YVXQNKPRZjIN4a9T93jjvrVddfqG8v3UZhREii++WIk7eISCAHa5F1U+uv4NydHCosTBMl7GA
QNKqcfBhb8K0hgR317uP89aBwxrNRCtQcVmGl3MPHGGWgjb3/utuhcVU4fng905gsh8Mo7xQOxJ5
S0VsVZXk6tIvc8X4pZMEwZ7PoGLwYSDAZAyqRkv0dlS0tv+9vGyzIPf0TsHJme5SljxOLkwYMf6N
60U4XOwJdb6GTUZ2u66NsDiSbm+T7vJFAMh4E/RSlB+wsNugTw91Zk6NQdQlzrBk5v5rAkck
`protect end_protected
