--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2014 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cc_cmplr_v3_0_7a1c77196b2a4f1a.vhd when simulating
-- the core, cc_cmplr_v3_0_7a1c77196b2a4f1a. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cc_cmplr_v3_0_7a1c77196b2a4f1a IS
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(87 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END cc_cmplr_v3_0_7a1c77196b2a4f1a;

ARCHITECTURE cc_cmplr_v3_0_7a1c77196b2a4f1a_a OF cc_cmplr_v3_0_7a1c77196b2a4f1a IS
-- synthesis translate_off
COMPONENT wrapped_cc_cmplr_v3_0_7a1c77196b2a4f1a
  PORT (
    aclk : IN STD_LOGIC;
    aclken : IN STD_LOGIC;
    s_axis_data_tdata : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
    s_axis_data_tvalid : IN STD_LOGIC;
    s_axis_data_tready : OUT STD_LOGIC;
    s_axis_data_tlast : IN STD_LOGIC;
    m_axis_data_tdata : OUT STD_LOGIC_VECTOR(87 DOWNTO 0);
    m_axis_data_tuser : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid : OUT STD_LOGIC;
    m_axis_data_tlast : OUT STD_LOGIC;
    event_tlast_unexpected : OUT STD_LOGIC;
    event_tlast_missing : OUT STD_LOGIC
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cc_cmplr_v3_0_7a1c77196b2a4f1a USE ENTITY XilinxCoreLib.cic_compiler_v3_0(behavioral)
    GENERIC MAP (
      c_c1 => 86,
      c_c2 => 86,
      c_c3 => 86,
      c_c4 => 86,
      c_c5 => 86,
      c_c6 => 0,
      c_clk_freq => 2000,
      c_component_name => "cc_cmplr_v3_0_7a1c77196b2a4f1a",
      c_diff_delay => 2,
      c_family => "virtex6",
      c_filter_type => 1,
      c_has_aclken => 1,
      c_has_aresetn => 0,
      c_has_dout_tready => 0,
      c_has_rounding => 0,
      c_i1 => 86,
      c_i2 => 86,
      c_i3 => 86,
      c_i4 => 86,
      c_i5 => 86,
      c_i6 => 0,
      c_input_width => 24,
      c_m_axis_data_tdata_width => 88,
      c_m_axis_data_tuser_width => 16,
      c_max_rate => 2500,
      c_min_rate => 2500,
      c_num_channels => 4,
      c_num_stages => 5,
      c_output_width => 86,
      c_rate => 2500,
      c_rate_type => 0,
      c_s_axis_config_tdata_width => 1,
      c_s_axis_data_tdata_width => 24,
      c_sample_freq => 1,
      c_use_dsp => 1,
      c_use_streaming_interface => 1,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cc_cmplr_v3_0_7a1c77196b2a4f1a
  PORT MAP (
    aclk => aclk,
    aclken => aclken,
    s_axis_data_tdata => s_axis_data_tdata,
    s_axis_data_tvalid => s_axis_data_tvalid,
    s_axis_data_tready => s_axis_data_tready,
    s_axis_data_tlast => s_axis_data_tlast,
    m_axis_data_tdata => m_axis_data_tdata,
    m_axis_data_tuser => m_axis_data_tuser,
    m_axis_data_tvalid => m_axis_data_tvalid,
    m_axis_data_tlast => m_axis_data_tlast,
    event_tlast_unexpected => event_tlast_unexpected,
    event_tlast_missing => event_tlast_missing
  );
-- synthesis translate_on

END cc_cmplr_v3_0_7a1c77196b2a4f1a_a;
