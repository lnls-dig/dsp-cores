`define ADDR_POS_CALC_DS_TBT_THRES     8'h0
`define POS_CALC_DS_TBT_THRES_VAL_OFFSET 0
`define POS_CALC_DS_TBT_THRES_VAL 32'h03ffffff
`define POS_CALC_DS_TBT_THRES_RESERVED_OFFSET 26
`define POS_CALC_DS_TBT_THRES_RESERVED 32'hfc000000
`define ADDR_POS_CALC_DS_FOFB_THRES    8'h4
`define POS_CALC_DS_FOFB_THRES_VAL_OFFSET 0
`define POS_CALC_DS_FOFB_THRES_VAL 32'h03ffffff
`define POS_CALC_DS_FOFB_THRES_RESERVED_OFFSET 26
`define POS_CALC_DS_FOFB_THRES_RESERVED 32'hfc000000
`define ADDR_POS_CALC_DS_MONIT_THRES   8'h8
`define POS_CALC_DS_MONIT_THRES_VAL_OFFSET 0
`define POS_CALC_DS_MONIT_THRES_VAL 32'h03ffffff
`define POS_CALC_DS_MONIT_THRES_RESERVED_OFFSET 26
`define POS_CALC_DS_MONIT_THRES_RESERVED 32'hfc000000
`define ADDR_POS_CALC_KX               8'hc
`define POS_CALC_KX_VAL_OFFSET 0
`define POS_CALC_KX_VAL 32'h01ffffff
`define POS_CALC_KX_RESERVED_OFFSET 25
`define POS_CALC_KX_RESERVED 32'hfe000000
`define ADDR_POS_CALC_KY               8'h10
`define POS_CALC_KY_VAL_OFFSET 0
`define POS_CALC_KY_VAL 32'h01ffffff
`define POS_CALC_KY_RESERVED_OFFSET 25
`define POS_CALC_KY_RESERVED 32'hfe000000
`define ADDR_POS_CALC_KSUM             8'h14
`define POS_CALC_KSUM_VAL_OFFSET 0
`define POS_CALC_KSUM_VAL 32'h01ffffff
`define POS_CALC_KSUM_RESERVED_OFFSET 25
`define POS_CALC_KSUM_RESERVED 32'hfe000000
`define ADDR_POS_CALC_DSP_CTNR_TBT     8'h18
`define POS_CALC_DSP_CTNR_TBT_CH01_OFFSET 0
`define POS_CALC_DSP_CTNR_TBT_CH01 32'h0000ffff
`define POS_CALC_DSP_CTNR_TBT_CH23_OFFSET 16
`define POS_CALC_DSP_CTNR_TBT_CH23 32'hffff0000
`define ADDR_POS_CALC_DSP_CTNR_FOFB    8'h1c
`define POS_CALC_DSP_CTNR_FOFB_CH01_OFFSET 0
`define POS_CALC_DSP_CTNR_FOFB_CH01 32'h0000ffff
`define POS_CALC_DSP_CTNR_FOFB_CH23_OFFSET 16
`define POS_CALC_DSP_CTNR_FOFB_CH23 32'hffff0000
`define ADDR_POS_CALC_DSP_CTNR1_MONIT  8'h20
`define POS_CALC_DSP_CTNR1_MONIT_CIC_OFFSET 0
`define POS_CALC_DSP_CTNR1_MONIT_CIC 32'h0000ffff
`define POS_CALC_DSP_CTNR1_MONIT_CFIR_OFFSET 16
`define POS_CALC_DSP_CTNR1_MONIT_CFIR 32'hffff0000
`define ADDR_POS_CALC_DSP_CTNR2_MONIT  8'h24
`define POS_CALC_DSP_CTNR2_MONIT_PFIR_OFFSET 0
`define POS_CALC_DSP_CTNR2_MONIT_PFIR 32'h0000ffff
`define POS_CALC_DSP_CTNR2_MONIT_FIR_01_OFFSET 16
`define POS_CALC_DSP_CTNR2_MONIT_FIR_01 32'hffff0000
`define ADDR_POS_CALC_DSP_ERR_CLR      8'h28
`define POS_CALC_DSP_ERR_CLR_TBT_OFFSET 0
`define POS_CALC_DSP_ERR_CLR_TBT 32'h00000001
`define POS_CALC_DSP_ERR_CLR_FOFB_OFFSET 1
`define POS_CALC_DSP_ERR_CLR_FOFB 32'h00000002
`define POS_CALC_DSP_ERR_CLR_MONIT_PART1_OFFSET 2
`define POS_CALC_DSP_ERR_CLR_MONIT_PART1 32'h00000004
`define POS_CALC_DSP_ERR_CLR_MONIT_PART2_OFFSET 3
`define POS_CALC_DSP_ERR_CLR_MONIT_PART2 32'h00000008
`define ADDR_POS_CALC_DDS_CFG          8'h2c
`define POS_CALC_DDS_CFG_VALID_CH0_OFFSET 0
`define POS_CALC_DDS_CFG_VALID_CH0 32'h00000001
`define POS_CALC_DDS_CFG_TEST_DATA_OFFSET 1
`define POS_CALC_DDS_CFG_TEST_DATA 32'h00000002
`define POS_CALC_DDS_CFG_RESERVED_CH0_OFFSET 2
`define POS_CALC_DDS_CFG_RESERVED_CH0 32'h000000fc
`define POS_CALC_DDS_CFG_VALID_CH1_OFFSET 8
`define POS_CALC_DDS_CFG_VALID_CH1 32'h00000100
`define POS_CALC_DDS_CFG_RESERVED_CH1_OFFSET 9
`define POS_CALC_DDS_CFG_RESERVED_CH1 32'h0000fe00
`define POS_CALC_DDS_CFG_VALID_CH2_OFFSET 16
`define POS_CALC_DDS_CFG_VALID_CH2 32'h00010000
`define POS_CALC_DDS_CFG_RESERVED_CH2_OFFSET 17
`define POS_CALC_DDS_CFG_RESERVED_CH2 32'h00fe0000
`define POS_CALC_DDS_CFG_VALID_CH3_OFFSET 24
`define POS_CALC_DDS_CFG_VALID_CH3 32'h01000000
`define POS_CALC_DDS_CFG_RESERVED_CH3_OFFSET 25
`define POS_CALC_DDS_CFG_RESERVED_CH3 32'hfe000000
`define ADDR_POS_CALC_DDS_PINC_CH0     8'h30
`define POS_CALC_DDS_PINC_CH0_VAL_OFFSET 0
`define POS_CALC_DDS_PINC_CH0_VAL 32'h3fffffff
`define POS_CALC_DDS_PINC_CH0_RESERVED_OFFSET 30
`define POS_CALC_DDS_PINC_CH0_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_PINC_CH1     8'h34
`define POS_CALC_DDS_PINC_CH1_VAL_OFFSET 0
`define POS_CALC_DDS_PINC_CH1_VAL 32'h3fffffff
`define POS_CALC_DDS_PINC_CH1_RESERVED_OFFSET 30
`define POS_CALC_DDS_PINC_CH1_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_PINC_CH2     8'h38
`define POS_CALC_DDS_PINC_CH2_VAL_OFFSET 0
`define POS_CALC_DDS_PINC_CH2_VAL 32'h3fffffff
`define POS_CALC_DDS_PINC_CH2_RESERVED_OFFSET 30
`define POS_CALC_DDS_PINC_CH2_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_PINC_CH3     8'h3c
`define POS_CALC_DDS_PINC_CH3_VAL_OFFSET 0
`define POS_CALC_DDS_PINC_CH3_VAL 32'h3fffffff
`define POS_CALC_DDS_PINC_CH3_RESERVED_OFFSET 30
`define POS_CALC_DDS_PINC_CH3_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_POFF_CH0     8'h40
`define POS_CALC_DDS_POFF_CH0_VAL_OFFSET 0
`define POS_CALC_DDS_POFF_CH0_VAL 32'h3fffffff
`define POS_CALC_DDS_POFF_CH0_RESERVED_OFFSET 30
`define POS_CALC_DDS_POFF_CH0_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_POFF_CH1     8'h44
`define POS_CALC_DDS_POFF_CH1_VAL_OFFSET 0
`define POS_CALC_DDS_POFF_CH1_VAL 32'h3fffffff
`define POS_CALC_DDS_POFF_CH1_RESERVED_OFFSET 30
`define POS_CALC_DDS_POFF_CH1_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_POFF_CH2     8'h48
`define POS_CALC_DDS_POFF_CH2_VAL_OFFSET 0
`define POS_CALC_DDS_POFF_CH2_VAL 32'h3fffffff
`define POS_CALC_DDS_POFF_CH2_RESERVED_OFFSET 30
`define POS_CALC_DDS_POFF_CH2_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DDS_POFF_CH3     8'h4c
`define POS_CALC_DDS_POFF_CH3_VAL_OFFSET 0
`define POS_CALC_DDS_POFF_CH3_VAL 32'h3fffffff
`define POS_CALC_DDS_POFF_CH3_RESERVED_OFFSET 30
`define POS_CALC_DDS_POFF_CH3_RESERVED 32'hc0000000
`define ADDR_POS_CALC_DSP_MONIT_AMP_CH0 8'h50
`define ADDR_POS_CALC_DSP_MONIT_AMP_CH1 8'h54
`define ADDR_POS_CALC_DSP_MONIT_AMP_CH2 8'h58
`define ADDR_POS_CALC_DSP_MONIT_AMP_CH3 8'h5c
`define ADDR_POS_CALC_DSP_MONIT_POS_X  8'h60
`define ADDR_POS_CALC_DSP_MONIT_POS_Y  8'h64
`define ADDR_POS_CALC_DSP_MONIT_POS_Q  8'h68
`define ADDR_POS_CALC_DSP_MONIT_POS_SUM 8'h6c
`define ADDR_POS_CALC_DSP_MONIT_UPDT   8'h70
`define ADDR_POS_CALC_DSP_MONIT1_AMP_CH0 8'h74
`define ADDR_POS_CALC_DSP_MONIT1_AMP_CH1 8'h78
`define ADDR_POS_CALC_DSP_MONIT1_AMP_CH2 8'h7c
`define ADDR_POS_CALC_DSP_MONIT1_AMP_CH3 8'h80
`define ADDR_POS_CALC_DSP_MONIT1_POS_X 8'h84
`define ADDR_POS_CALC_DSP_MONIT1_POS_Y 8'h88
`define ADDR_POS_CALC_DSP_MONIT1_POS_Q 8'h8c
`define ADDR_POS_CALC_DSP_MONIT1_POS_SUM 8'h90
`define ADDR_POS_CALC_DSP_MONIT1_UPDT  8'h94
`define ADDR_POS_CALC_AMPFIFO_MONIT_R0 8'h98
`define POS_CALC_AMPFIFO_MONIT_R0_AMP_CH0_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT_R0_AMP_CH0 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT_R1 8'h9c
`define POS_CALC_AMPFIFO_MONIT_R1_AMP_CH1_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT_R1_AMP_CH1 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT_R2 8'ha0
`define POS_CALC_AMPFIFO_MONIT_R2_AMP_CH2_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT_R2_AMP_CH2 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT_R3 8'ha4
`define POS_CALC_AMPFIFO_MONIT_R3_AMP_CH3_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT_R3_AMP_CH3 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT_CSR 8'ha8
`define POS_CALC_AMPFIFO_MONIT_CSR_FULL_OFFSET 16
`define POS_CALC_AMPFIFO_MONIT_CSR_FULL 32'h00010000
`define POS_CALC_AMPFIFO_MONIT_CSR_EMPTY_OFFSET 17
`define POS_CALC_AMPFIFO_MONIT_CSR_EMPTY 32'h00020000
`define POS_CALC_AMPFIFO_MONIT_CSR_USEDW_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT_CSR_USEDW 32'h0000000f
`define ADDR_POS_CALC_POSFIFO_MONIT_R0 8'hac
`define POS_CALC_POSFIFO_MONIT_R0_POS_X_OFFSET 0
`define POS_CALC_POSFIFO_MONIT_R0_POS_X 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT_R1 8'hb0
`define POS_CALC_POSFIFO_MONIT_R1_POS_Y_OFFSET 0
`define POS_CALC_POSFIFO_MONIT_R1_POS_Y 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT_R2 8'hb4
`define POS_CALC_POSFIFO_MONIT_R2_POS_Q_OFFSET 0
`define POS_CALC_POSFIFO_MONIT_R2_POS_Q 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT_R3 8'hb8
`define POS_CALC_POSFIFO_MONIT_R3_POS_SUM_OFFSET 0
`define POS_CALC_POSFIFO_MONIT_R3_POS_SUM 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT_CSR 8'hbc
`define POS_CALC_POSFIFO_MONIT_CSR_FULL_OFFSET 16
`define POS_CALC_POSFIFO_MONIT_CSR_FULL 32'h00010000
`define POS_CALC_POSFIFO_MONIT_CSR_EMPTY_OFFSET 17
`define POS_CALC_POSFIFO_MONIT_CSR_EMPTY 32'h00020000
`define POS_CALC_POSFIFO_MONIT_CSR_USEDW_OFFSET 0
`define POS_CALC_POSFIFO_MONIT_CSR_USEDW 32'h0000000f
`define ADDR_POS_CALC_AMPFIFO_MONIT1_R0 8'hc0
`define POS_CALC_AMPFIFO_MONIT1_R0_AMP_CH0_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT1_R0_AMP_CH0 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT1_R1 8'hc4
`define POS_CALC_AMPFIFO_MONIT1_R1_AMP_CH1_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT1_R1_AMP_CH1 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT1_R2 8'hc8
`define POS_CALC_AMPFIFO_MONIT1_R2_AMP_CH2_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT1_R2_AMP_CH2 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT1_R3 8'hcc
`define POS_CALC_AMPFIFO_MONIT1_R3_AMP_CH3_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT1_R3_AMP_CH3 32'hffffffff
`define ADDR_POS_CALC_AMPFIFO_MONIT1_CSR 8'hd0
`define POS_CALC_AMPFIFO_MONIT1_CSR_FULL_OFFSET 16
`define POS_CALC_AMPFIFO_MONIT1_CSR_FULL 32'h00010000
`define POS_CALC_AMPFIFO_MONIT1_CSR_EMPTY_OFFSET 17
`define POS_CALC_AMPFIFO_MONIT1_CSR_EMPTY 32'h00020000
`define POS_CALC_AMPFIFO_MONIT1_CSR_USEDW_OFFSET 0
`define POS_CALC_AMPFIFO_MONIT1_CSR_USEDW 32'h0000000f
`define ADDR_POS_CALC_POSFIFO_MONIT1_R0 8'hd4
`define POS_CALC_POSFIFO_MONIT1_R0_POS_X_OFFSET 0
`define POS_CALC_POSFIFO_MONIT1_R0_POS_X 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT1_R1 8'hd8
`define POS_CALC_POSFIFO_MONIT1_R1_POS_Y_OFFSET 0
`define POS_CALC_POSFIFO_MONIT1_R1_POS_Y 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT1_R2 8'hdc
`define POS_CALC_POSFIFO_MONIT1_R2_POS_Q_OFFSET 0
`define POS_CALC_POSFIFO_MONIT1_R2_POS_Q 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT1_R3 8'he0
`define POS_CALC_POSFIFO_MONIT1_R3_POS_SUM_OFFSET 0
`define POS_CALC_POSFIFO_MONIT1_R3_POS_SUM 32'hffffffff
`define ADDR_POS_CALC_POSFIFO_MONIT1_CSR 8'he4
`define POS_CALC_POSFIFO_MONIT1_CSR_FULL_OFFSET 16
`define POS_CALC_POSFIFO_MONIT1_CSR_FULL 32'h00010000
`define POS_CALC_POSFIFO_MONIT1_CSR_EMPTY_OFFSET 17
`define POS_CALC_POSFIFO_MONIT1_CSR_EMPTY 32'h00020000
`define POS_CALC_POSFIFO_MONIT1_CSR_USEDW_OFFSET 0
`define POS_CALC_POSFIFO_MONIT1_CSR_USEDW 32'h0000000f
`define ADDR_POS_CALC_SW_TAG           8'he8
`define POS_CALC_SW_TAG_EN_OFFSET 0
`define POS_CALC_SW_TAG_EN 32'h00000001
`define POS_CALC_SW_TAG_DESYNC_CNT_RST_OFFSET 8
`define POS_CALC_SW_TAG_DESYNC_CNT_RST 32'h00000100
`define POS_CALC_SW_TAG_DESYNC_CNT_OFFSET 9
`define POS_CALC_SW_TAG_DESYNC_CNT 32'h007ffe00
`define ADDR_POS_CALC_SW_DATA_MASK     8'hec
`define POS_CALC_SW_DATA_MASK_EN_OFFSET 0
`define POS_CALC_SW_DATA_MASK_EN 32'h00000001
`define POS_CALC_SW_DATA_MASK_SAMPLES_OFFSET 1
`define POS_CALC_SW_DATA_MASK_SAMPLES 32'h0001fffe
`define ADDR_POS_CALC_TBT_TAG    8'hf0
`define POS_CALC_TBT_TAG_EN_OFFSET 0
`define POS_CALC_TBT_TAG_EN 32'h00000001
`define POS_CALC_TBT_TAG_DLY_OFFSET 1
`define POS_CALC_TBT_TAG_DLY 32'h0001fffe
`define POS_CALC_TBT_TAG_DESYNC_CNT_RST_OFFSET 17
`define POS_CALC_TBT_TAG_DESYNC_CNT_RST 32'h00020000
`define POS_CALC_TBT_TAG_DESYNC_CNT_OFFSET 18
`define POS_CALC_TBT_TAG_DESYNC_CNT 32'hfffc0000
`define ADDR_POS_CALC_TBT_DATA_MASK_CTL 8'hf4
`define POS_CALC_TBT_DATA_MASK_CTL_EN_OFFSET 0
`define POS_CALC_TBT_DATA_MASK_CTL_EN 32'h00000001
`define ADDR_POS_CALC_TBT_DATA_MASK_SAMPLES 8'hf8
`define POS_CALC_TBT_DATA_MASK_SAMPLES_BEG_OFFSET 0
`define POS_CALC_TBT_DATA_MASK_SAMPLES_BEG 32'h0000ffff
`define POS_CALC_TBT_DATA_MASK_SAMPLES_END_OFFSET 16
`define POS_CALC_TBT_DATA_MASK_SAMPLES_END 32'hffff0000
