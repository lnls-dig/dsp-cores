`define ADDR_BPM_SWAP_CTRL             5'h0
`define BPM_SWAP_CTRL_RST_OFFSET 0
`define BPM_SWAP_CTRL_RST 32'h00000001
`define BPM_SWAP_CTRL_MODE1_OFFSET 1
`define BPM_SWAP_CTRL_MODE1 32'h00000006
`define BPM_SWAP_CTRL_MODE2_OFFSET 3
`define BPM_SWAP_CTRL_MODE2 32'h00000018
`define BPM_SWAP_CTRL_SWAP_DIV_F_OFFSET 8
`define BPM_SWAP_CTRL_SWAP_DIV_F 32'h00ffff00
`define ADDR_BPM_SWAP_DLY              5'h4
`define BPM_SWAP_DLY_1_OFFSET 0
`define BPM_SWAP_DLY_1 32'h0000ffff
`define BPM_SWAP_DLY_2_OFFSET 16
`define BPM_SWAP_DLY_2 32'hffff0000
`define ADDR_BPM_SWAP_A                5'h8
`define BPM_SWAP_A_A_OFFSET 0
`define BPM_SWAP_A_A 32'h000003ff
`define BPM_SWAP_A_C_OFFSET 16
`define BPM_SWAP_A_C 32'h03ff0000
`define ADDR_BPM_SWAP_B                5'hc
`define BPM_SWAP_B_B_OFFSET 0
`define BPM_SWAP_B_B 32'h000003ff
`define BPM_SWAP_B_D_OFFSET 16
`define BPM_SWAP_B_D 32'h03ff0000
`define ADDR_BPM_SWAP_C                5'h10
`define BPM_SWAP_C_C_OFFSET 0
`define BPM_SWAP_C_C 32'h000003ff
`define BPM_SWAP_C_A_OFFSET 16
`define BPM_SWAP_C_A 32'h03ff0000
`define ADDR_BPM_SWAP_D                5'h14
`define BPM_SWAP_D_D_OFFSET 0
`define BPM_SWAP_D_D 32'h000003ff
`define BPM_SWAP_D_B_OFFSET 16
`define BPM_SWAP_D_B 32'h03ff0000
`define ADDR_BPM_SWAP_DUMMY            5'h18
